##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 23:52:37 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16_64
  CLASS BLOCK ;
  SIZE 154.6000 BY 86.6000 ;
  FOREIGN sram_w16_64 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 35.3500 0.6000 35.4500 ;
    END
  END CLK
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.8500 0.0000 125.9500 0.6000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.2500 0.0000 124.3500 0.6000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.6500 0.0000 122.7500 0.6000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.0500 0.0000 121.1500 0.6000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.4500 0.0000 119.5500 0.6000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.8500 0.0000 117.9500 0.6000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.2500 0.0000 116.3500 0.6000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.6500 0.0000 114.7500 0.6000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.0500 0.0000 113.1500 0.6000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.4500 0.0000 111.5500 0.6000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.8500 0.0000 109.9500 0.6000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.2500 0.0000 108.3500 0.6000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.6500 0.0000 106.7500 0.6000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.0500 0.0000 105.1500 0.6000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.4500 0.0000 103.5500 0.6000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.8500 0.0000 101.9500 0.6000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.2500 0.0000 100.3500 0.6000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.6500 0.0000 98.7500 0.6000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.0500 0.0000 97.1500 0.6000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.4500 0.0000 95.5500 0.6000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.8500 0.0000 93.9500 0.6000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.2500 0.0000 92.3500 0.6000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.6500 0.0000 90.7500 0.6000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.0500 0.0000 89.1500 0.6000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.4500 0.0000 87.5500 0.6000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.8500 0.0000 85.9500 0.6000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.2500 0.0000 84.3500 0.6000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.6500 0.0000 82.7500 0.6000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.0500 0.0000 81.1500 0.6000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.4500 0.0000 79.5500 0.6000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 77.8500 0.0000 77.9500 0.6000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.2500 0.0000 76.3500 0.6000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 74.6500 0.0000 74.7500 0.6000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.0500 0.0000 73.1500 0.6000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.4500 0.0000 71.5500 0.6000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 69.8500 0.0000 69.9500 0.6000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.2500 0.0000 68.3500 0.6000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 66.6500 0.0000 66.7500 0.6000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.0500 0.0000 65.1500 0.6000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 63.4500 0.0000 63.5500 0.6000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 61.8500 0.0000 61.9500 0.6000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60.2500 0.0000 60.3500 0.6000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.6500 0.0000 58.7500 0.6000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 57.0500 0.0000 57.1500 0.6000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.4500 0.0000 55.5500 0.6000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 53.8500 0.0000 53.9500 0.6000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.2500 0.0000 52.3500 0.6000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 50.6500 0.0000 50.7500 0.6000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 49.0500 0.0000 49.1500 0.6000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 47.4500 0.0000 47.5500 0.6000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 45.8500 0.0000 45.9500 0.6000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 44.2500 0.0000 44.3500 0.6000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 42.6500 0.0000 42.7500 0.6000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 41.0500 0.0000 41.1500 0.6000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.4500 0.0000 39.5500 0.6000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 37.8500 0.0000 37.9500 0.6000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 36.2500 0.0000 36.3500 0.6000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 34.6500 0.0000 34.7500 0.6000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 33.0500 0.0000 33.1500 0.6000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 31.4500 0.0000 31.5500 0.6000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 29.8500 0.0000 29.9500 0.6000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 28.2500 0.0000 28.3500 0.6000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 26.6500 0.0000 26.7500 0.6000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 25.0500 0.0000 25.1500 0.6000 ;
    END
  END D[0]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.8500 86.0000 125.9500 86.6000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.2500 86.0000 124.3500 86.6000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.6500 86.0000 122.7500 86.6000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.0500 86.0000 121.1500 86.6000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.4500 86.0000 119.5500 86.6000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.8500 86.0000 117.9500 86.6000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.2500 86.0000 116.3500 86.6000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.6500 86.0000 114.7500 86.6000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.0500 86.0000 113.1500 86.6000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.4500 86.0000 111.5500 86.6000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.8500 86.0000 109.9500 86.6000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.2500 86.0000 108.3500 86.6000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.6500 86.0000 106.7500 86.6000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.0500 86.0000 105.1500 86.6000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.4500 86.0000 103.5500 86.6000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.8500 86.0000 101.9500 86.6000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.2500 86.0000 100.3500 86.6000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.6500 86.0000 98.7500 86.6000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.0500 86.0000 97.1500 86.6000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.4500 86.0000 95.5500 86.6000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.8500 86.0000 93.9500 86.6000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.2500 86.0000 92.3500 86.6000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.6500 86.0000 90.7500 86.6000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.0500 86.0000 89.1500 86.6000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.4500 86.0000 87.5500 86.6000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.8500 86.0000 85.9500 86.6000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.2500 86.0000 84.3500 86.6000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.6500 86.0000 82.7500 86.6000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.0500 86.0000 81.1500 86.6000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.4500 86.0000 79.5500 86.6000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 77.8500 86.0000 77.9500 86.6000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.2500 86.0000 76.3500 86.6000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 74.6500 86.0000 74.7500 86.6000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.0500 86.0000 73.1500 86.6000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.4500 86.0000 71.5500 86.6000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 69.8500 86.0000 69.9500 86.6000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.2500 86.0000 68.3500 86.6000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 66.6500 86.0000 66.7500 86.6000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.0500 86.0000 65.1500 86.6000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 63.4500 86.0000 63.5500 86.6000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 61.8500 86.0000 61.9500 86.6000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60.2500 86.0000 60.3500 86.6000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.6500 86.0000 58.7500 86.6000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 57.0500 86.0000 57.1500 86.6000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.4500 86.0000 55.5500 86.6000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 53.8500 86.0000 53.9500 86.6000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.2500 86.0000 52.3500 86.6000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 50.6500 86.0000 50.7500 86.6000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 49.0500 86.0000 49.1500 86.6000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 47.4500 86.0000 47.5500 86.6000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 45.8500 86.0000 45.9500 86.6000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 44.2500 86.0000 44.3500 86.6000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 42.6500 86.0000 42.7500 86.6000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 41.0500 86.0000 41.1500 86.6000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.4500 86.0000 39.5500 86.6000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 37.8500 86.0000 37.9500 86.6000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 36.2500 86.0000 36.3500 86.6000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 34.6500 86.0000 34.7500 86.6000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 33.0500 86.0000 33.1500 86.6000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 31.4500 86.0000 31.5500 86.6000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 29.8500 86.0000 29.9500 86.6000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 28.2500 86.0000 28.3500 86.6000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 26.6500 86.0000 26.7500 86.6000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 25.0500 86.0000 25.1500 86.6000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 39.3500 0.6000 39.4500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.3500 0.6000 31.4500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 43.3500 0.6000 43.4500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 47.3500 0.6000 47.4500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 51.3500 0.6000 51.4500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.3500 0.6000 55.4500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 30.0000 10.0000 32.0000 76.6000 ;
        RECT 58.5300 10.0000 60.5300 76.6000 ;
        RECT 87.0600 10.0000 89.0600 76.6000 ;
        RECT 115.5900 10.0000 117.5900 76.6000 ;
        RECT 30.0000 76.4350 32.0000 76.7650 ;
        RECT 58.5300 76.4350 60.5300 76.7650 ;
        RECT 115.5900 76.4350 117.5900 76.7650 ;
        RECT 87.0600 76.4350 89.0600 76.7650 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 37.0000 10.0000 39.0000 76.6000 ;
        RECT 65.5300 10.0000 67.5300 76.6000 ;
        RECT 94.0600 10.0000 96.0600 76.6000 ;
        RECT 122.5900 10.0000 124.5900 76.6000 ;
        RECT 37.0000 9.8350 39.0000 10.1650 ;
        RECT 65.5300 9.8350 67.5300 10.1650 ;
        RECT 94.0600 9.8350 96.0600 10.1650 ;
        RECT 122.5900 9.8350 124.5900 10.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 154.6000 86.6000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 154.6000 86.6000 ;
    LAYER M3 ;
      RECT 126.1100 85.8400 154.6000 86.6000 ;
      RECT 124.5100 85.8400 125.6900 86.6000 ;
      RECT 122.9100 85.8400 124.0900 86.6000 ;
      RECT 121.3100 85.8400 122.4900 86.6000 ;
      RECT 119.7100 85.8400 120.8900 86.6000 ;
      RECT 118.1100 85.8400 119.2900 86.6000 ;
      RECT 116.5100 85.8400 117.6900 86.6000 ;
      RECT 114.9100 85.8400 116.0900 86.6000 ;
      RECT 113.3100 85.8400 114.4900 86.6000 ;
      RECT 111.7100 85.8400 112.8900 86.6000 ;
      RECT 110.1100 85.8400 111.2900 86.6000 ;
      RECT 108.5100 85.8400 109.6900 86.6000 ;
      RECT 106.9100 85.8400 108.0900 86.6000 ;
      RECT 105.3100 85.8400 106.4900 86.6000 ;
      RECT 103.7100 85.8400 104.8900 86.6000 ;
      RECT 102.1100 85.8400 103.2900 86.6000 ;
      RECT 100.5100 85.8400 101.6900 86.6000 ;
      RECT 98.9100 85.8400 100.0900 86.6000 ;
      RECT 97.3100 85.8400 98.4900 86.6000 ;
      RECT 95.7100 85.8400 96.8900 86.6000 ;
      RECT 94.1100 85.8400 95.2900 86.6000 ;
      RECT 92.5100 85.8400 93.6900 86.6000 ;
      RECT 90.9100 85.8400 92.0900 86.6000 ;
      RECT 89.3100 85.8400 90.4900 86.6000 ;
      RECT 87.7100 85.8400 88.8900 86.6000 ;
      RECT 86.1100 85.8400 87.2900 86.6000 ;
      RECT 84.5100 85.8400 85.6900 86.6000 ;
      RECT 82.9100 85.8400 84.0900 86.6000 ;
      RECT 81.3100 85.8400 82.4900 86.6000 ;
      RECT 79.7100 85.8400 80.8900 86.6000 ;
      RECT 78.1100 85.8400 79.2900 86.6000 ;
      RECT 76.5100 85.8400 77.6900 86.6000 ;
      RECT 74.9100 85.8400 76.0900 86.6000 ;
      RECT 73.3100 85.8400 74.4900 86.6000 ;
      RECT 71.7100 85.8400 72.8900 86.6000 ;
      RECT 70.1100 85.8400 71.2900 86.6000 ;
      RECT 68.5100 85.8400 69.6900 86.6000 ;
      RECT 66.9100 85.8400 68.0900 86.6000 ;
      RECT 65.3100 85.8400 66.4900 86.6000 ;
      RECT 63.7100 85.8400 64.8900 86.6000 ;
      RECT 62.1100 85.8400 63.2900 86.6000 ;
      RECT 60.5100 85.8400 61.6900 86.6000 ;
      RECT 58.9100 85.8400 60.0900 86.6000 ;
      RECT 57.3100 85.8400 58.4900 86.6000 ;
      RECT 55.7100 85.8400 56.8900 86.6000 ;
      RECT 54.1100 85.8400 55.2900 86.6000 ;
      RECT 52.5100 85.8400 53.6900 86.6000 ;
      RECT 50.9100 85.8400 52.0900 86.6000 ;
      RECT 49.3100 85.8400 50.4900 86.6000 ;
      RECT 47.7100 85.8400 48.8900 86.6000 ;
      RECT 46.1100 85.8400 47.2900 86.6000 ;
      RECT 44.5100 85.8400 45.6900 86.6000 ;
      RECT 42.9100 85.8400 44.0900 86.6000 ;
      RECT 41.3100 85.8400 42.4900 86.6000 ;
      RECT 39.7100 85.8400 40.8900 86.6000 ;
      RECT 38.1100 85.8400 39.2900 86.6000 ;
      RECT 36.5100 85.8400 37.6900 86.6000 ;
      RECT 34.9100 85.8400 36.0900 86.6000 ;
      RECT 33.3100 85.8400 34.4900 86.6000 ;
      RECT 31.7100 85.8400 32.8900 86.6000 ;
      RECT 30.1100 85.8400 31.2900 86.6000 ;
      RECT 28.5100 85.8400 29.6900 86.6000 ;
      RECT 26.9100 85.8400 28.0900 86.6000 ;
      RECT 25.3100 85.8400 26.4900 86.6000 ;
      RECT 0.0000 85.8400 24.8900 86.6000 ;
      RECT 0.0000 55.5500 154.6000 85.8400 ;
      RECT 0.7000 55.2500 154.6000 55.5500 ;
      RECT 0.0000 51.5500 154.6000 55.2500 ;
      RECT 0.7000 51.2500 154.6000 51.5500 ;
      RECT 0.0000 47.5500 154.6000 51.2500 ;
      RECT 0.7000 47.2500 154.6000 47.5500 ;
      RECT 0.0000 43.5500 154.6000 47.2500 ;
      RECT 0.7000 43.2500 154.6000 43.5500 ;
      RECT 0.0000 39.5500 154.6000 43.2500 ;
      RECT 0.7000 39.2500 154.6000 39.5500 ;
      RECT 0.0000 35.5500 154.6000 39.2500 ;
      RECT 0.7000 35.2500 154.6000 35.5500 ;
      RECT 0.0000 31.5500 154.6000 35.2500 ;
      RECT 0.7000 31.2500 154.6000 31.5500 ;
      RECT 0.0000 0.7600 154.6000 31.2500 ;
      RECT 126.1100 0.0000 154.6000 0.7600 ;
      RECT 124.5100 0.0000 125.6900 0.7600 ;
      RECT 122.9100 0.0000 124.0900 0.7600 ;
      RECT 121.3100 0.0000 122.4900 0.7600 ;
      RECT 119.7100 0.0000 120.8900 0.7600 ;
      RECT 118.1100 0.0000 119.2900 0.7600 ;
      RECT 116.5100 0.0000 117.6900 0.7600 ;
      RECT 114.9100 0.0000 116.0900 0.7600 ;
      RECT 113.3100 0.0000 114.4900 0.7600 ;
      RECT 111.7100 0.0000 112.8900 0.7600 ;
      RECT 110.1100 0.0000 111.2900 0.7600 ;
      RECT 108.5100 0.0000 109.6900 0.7600 ;
      RECT 106.9100 0.0000 108.0900 0.7600 ;
      RECT 105.3100 0.0000 106.4900 0.7600 ;
      RECT 103.7100 0.0000 104.8900 0.7600 ;
      RECT 102.1100 0.0000 103.2900 0.7600 ;
      RECT 100.5100 0.0000 101.6900 0.7600 ;
      RECT 98.9100 0.0000 100.0900 0.7600 ;
      RECT 97.3100 0.0000 98.4900 0.7600 ;
      RECT 95.7100 0.0000 96.8900 0.7600 ;
      RECT 94.1100 0.0000 95.2900 0.7600 ;
      RECT 92.5100 0.0000 93.6900 0.7600 ;
      RECT 90.9100 0.0000 92.0900 0.7600 ;
      RECT 89.3100 0.0000 90.4900 0.7600 ;
      RECT 87.7100 0.0000 88.8900 0.7600 ;
      RECT 86.1100 0.0000 87.2900 0.7600 ;
      RECT 84.5100 0.0000 85.6900 0.7600 ;
      RECT 82.9100 0.0000 84.0900 0.7600 ;
      RECT 81.3100 0.0000 82.4900 0.7600 ;
      RECT 79.7100 0.0000 80.8900 0.7600 ;
      RECT 78.1100 0.0000 79.2900 0.7600 ;
      RECT 76.5100 0.0000 77.6900 0.7600 ;
      RECT 74.9100 0.0000 76.0900 0.7600 ;
      RECT 73.3100 0.0000 74.4900 0.7600 ;
      RECT 71.7100 0.0000 72.8900 0.7600 ;
      RECT 70.1100 0.0000 71.2900 0.7600 ;
      RECT 68.5100 0.0000 69.6900 0.7600 ;
      RECT 66.9100 0.0000 68.0900 0.7600 ;
      RECT 65.3100 0.0000 66.4900 0.7600 ;
      RECT 63.7100 0.0000 64.8900 0.7600 ;
      RECT 62.1100 0.0000 63.2900 0.7600 ;
      RECT 60.5100 0.0000 61.6900 0.7600 ;
      RECT 58.9100 0.0000 60.0900 0.7600 ;
      RECT 57.3100 0.0000 58.4900 0.7600 ;
      RECT 55.7100 0.0000 56.8900 0.7600 ;
      RECT 54.1100 0.0000 55.2900 0.7600 ;
      RECT 52.5100 0.0000 53.6900 0.7600 ;
      RECT 50.9100 0.0000 52.0900 0.7600 ;
      RECT 49.3100 0.0000 50.4900 0.7600 ;
      RECT 47.7100 0.0000 48.8900 0.7600 ;
      RECT 46.1100 0.0000 47.2900 0.7600 ;
      RECT 44.5100 0.0000 45.6900 0.7600 ;
      RECT 42.9100 0.0000 44.0900 0.7600 ;
      RECT 41.3100 0.0000 42.4900 0.7600 ;
      RECT 39.7100 0.0000 40.8900 0.7600 ;
      RECT 38.1100 0.0000 39.2900 0.7600 ;
      RECT 36.5100 0.0000 37.6900 0.7600 ;
      RECT 34.9100 0.0000 36.0900 0.7600 ;
      RECT 33.3100 0.0000 34.4900 0.7600 ;
      RECT 31.7100 0.0000 32.8900 0.7600 ;
      RECT 30.1100 0.0000 31.2900 0.7600 ;
      RECT 28.5100 0.0000 29.6900 0.7600 ;
      RECT 26.9100 0.0000 28.0900 0.7600 ;
      RECT 25.3100 0.0000 26.4900 0.7600 ;
      RECT 0.0000 0.0000 24.8900 0.7600 ;
    LAYER M4 ;
      RECT 0.0000 77.2650 154.6000 86.6000 ;
      RECT 118.0900 77.1000 154.6000 77.2650 ;
      RECT 89.5600 77.1000 115.0900 77.2650 ;
      RECT 61.0300 77.1000 86.5600 77.2650 ;
      RECT 32.5000 77.1000 58.0300 77.2650 ;
      RECT 118.0900 9.5000 122.0900 77.1000 ;
      RECT 96.5600 9.5000 115.0900 77.1000 ;
      RECT 89.5600 9.5000 93.5600 77.1000 ;
      RECT 68.0300 9.5000 86.5600 77.1000 ;
      RECT 61.0300 9.5000 65.0300 77.1000 ;
      RECT 39.5000 9.5000 58.0300 77.1000 ;
      RECT 32.5000 9.5000 36.5000 77.1000 ;
      RECT 0.0000 9.5000 29.5000 77.2650 ;
      RECT 125.0900 9.3350 154.6000 77.1000 ;
      RECT 96.5600 9.3350 122.0900 9.5000 ;
      RECT 68.0300 9.3350 93.5600 9.5000 ;
      RECT 39.5000 9.3350 65.0300 9.5000 ;
      RECT 0.0000 9.3350 36.5000 9.5000 ;
      RECT 0.0000 0.0000 154.6000 9.3350 ;
  END
END sram_w16_64

END LIBRARY
