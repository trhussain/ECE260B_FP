##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 19:10:39 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16_256
  CLASS BLOCK ;
  SIZE 450.2000 BY 102.8000 ;
  FOREIGN sram_w16_256 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 43.5500 0.6000 43.6500 ;
    END
  END CLK
  PIN D[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 433.0500 0.0000 433.1500 0.6000 ;
    END
  END D[255]
  PIN D[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 431.4500 0.0000 431.5500 0.6000 ;
    END
  END D[254]
  PIN D[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 429.8500 0.0000 429.9500 0.6000 ;
    END
  END D[253]
  PIN D[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 428.2500 0.0000 428.3500 0.6000 ;
    END
  END D[252]
  PIN D[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 426.6500 0.0000 426.7500 0.6000 ;
    END
  END D[251]
  PIN D[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 425.0500 0.0000 425.1500 0.6000 ;
    END
  END D[250]
  PIN D[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 423.4500 0.0000 423.5500 0.6000 ;
    END
  END D[249]
  PIN D[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 421.8500 0.0000 421.9500 0.6000 ;
    END
  END D[248]
  PIN D[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 420.2500 0.0000 420.3500 0.6000 ;
    END
  END D[247]
  PIN D[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 418.6500 0.0000 418.7500 0.6000 ;
    END
  END D[246]
  PIN D[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 417.0500 0.0000 417.1500 0.6000 ;
    END
  END D[245]
  PIN D[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 415.4500 0.0000 415.5500 0.6000 ;
    END
  END D[244]
  PIN D[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 413.8500 0.0000 413.9500 0.6000 ;
    END
  END D[243]
  PIN D[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 412.2500 0.0000 412.3500 0.6000 ;
    END
  END D[242]
  PIN D[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 410.6500 0.0000 410.7500 0.6000 ;
    END
  END D[241]
  PIN D[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 409.0500 0.0000 409.1500 0.6000 ;
    END
  END D[240]
  PIN D[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 407.4500 0.0000 407.5500 0.6000 ;
    END
  END D[239]
  PIN D[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 405.8500 0.0000 405.9500 0.6000 ;
    END
  END D[238]
  PIN D[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 404.2500 0.0000 404.3500 0.6000 ;
    END
  END D[237]
  PIN D[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 402.6500 0.0000 402.7500 0.6000 ;
    END
  END D[236]
  PIN D[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.0500 0.0000 401.1500 0.6000 ;
    END
  END D[235]
  PIN D[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 399.4500 0.0000 399.5500 0.6000 ;
    END
  END D[234]
  PIN D[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 397.8500 0.0000 397.9500 0.6000 ;
    END
  END D[233]
  PIN D[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 396.2500 0.0000 396.3500 0.6000 ;
    END
  END D[232]
  PIN D[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 394.6500 0.0000 394.7500 0.6000 ;
    END
  END D[231]
  PIN D[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 393.0500 0.0000 393.1500 0.6000 ;
    END
  END D[230]
  PIN D[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 391.4500 0.0000 391.5500 0.6000 ;
    END
  END D[229]
  PIN D[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 389.8500 0.0000 389.9500 0.6000 ;
    END
  END D[228]
  PIN D[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 388.2500 0.0000 388.3500 0.6000 ;
    END
  END D[227]
  PIN D[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 386.6500 0.0000 386.7500 0.6000 ;
    END
  END D[226]
  PIN D[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 385.0500 0.0000 385.1500 0.6000 ;
    END
  END D[225]
  PIN D[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 383.4500 0.0000 383.5500 0.6000 ;
    END
  END D[224]
  PIN D[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 381.8500 0.0000 381.9500 0.6000 ;
    END
  END D[223]
  PIN D[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380.2500 0.0000 380.3500 0.6000 ;
    END
  END D[222]
  PIN D[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 378.6500 0.0000 378.7500 0.6000 ;
    END
  END D[221]
  PIN D[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 377.0500 0.0000 377.1500 0.6000 ;
    END
  END D[220]
  PIN D[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 375.4500 0.0000 375.5500 0.6000 ;
    END
  END D[219]
  PIN D[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 373.8500 0.0000 373.9500 0.6000 ;
    END
  END D[218]
  PIN D[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 372.2500 0.0000 372.3500 0.6000 ;
    END
  END D[217]
  PIN D[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 370.6500 0.0000 370.7500 0.6000 ;
    END
  END D[216]
  PIN D[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 369.0500 0.0000 369.1500 0.6000 ;
    END
  END D[215]
  PIN D[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 367.4500 0.0000 367.5500 0.6000 ;
    END
  END D[214]
  PIN D[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 365.8500 0.0000 365.9500 0.6000 ;
    END
  END D[213]
  PIN D[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 364.2500 0.0000 364.3500 0.6000 ;
    END
  END D[212]
  PIN D[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 362.6500 0.0000 362.7500 0.6000 ;
    END
  END D[211]
  PIN D[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 361.0500 0.0000 361.1500 0.6000 ;
    END
  END D[210]
  PIN D[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 359.4500 0.0000 359.5500 0.6000 ;
    END
  END D[209]
  PIN D[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 357.8500 0.0000 357.9500 0.6000 ;
    END
  END D[208]
  PIN D[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 356.2500 0.0000 356.3500 0.6000 ;
    END
  END D[207]
  PIN D[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 354.6500 0.0000 354.7500 0.6000 ;
    END
  END D[206]
  PIN D[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 353.0500 0.0000 353.1500 0.6000 ;
    END
  END D[205]
  PIN D[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 351.4500 0.0000 351.5500 0.6000 ;
    END
  END D[204]
  PIN D[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 349.8500 0.0000 349.9500 0.6000 ;
    END
  END D[203]
  PIN D[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 348.2500 0.0000 348.3500 0.6000 ;
    END
  END D[202]
  PIN D[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 346.6500 0.0000 346.7500 0.6000 ;
    END
  END D[201]
  PIN D[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 345.0500 0.0000 345.1500 0.6000 ;
    END
  END D[200]
  PIN D[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 343.4500 0.0000 343.5500 0.6000 ;
    END
  END D[199]
  PIN D[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 341.8500 0.0000 341.9500 0.6000 ;
    END
  END D[198]
  PIN D[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 340.2500 0.0000 340.3500 0.6000 ;
    END
  END D[197]
  PIN D[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 338.6500 0.0000 338.7500 0.6000 ;
    END
  END D[196]
  PIN D[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 337.0500 0.0000 337.1500 0.6000 ;
    END
  END D[195]
  PIN D[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 335.4500 0.0000 335.5500 0.6000 ;
    END
  END D[194]
  PIN D[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 333.8500 0.0000 333.9500 0.6000 ;
    END
  END D[193]
  PIN D[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 332.2500 0.0000 332.3500 0.6000 ;
    END
  END D[192]
  PIN D[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 330.6500 0.0000 330.7500 0.6000 ;
    END
  END D[191]
  PIN D[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 329.0500 0.0000 329.1500 0.6000 ;
    END
  END D[190]
  PIN D[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.4500 0.0000 327.5500 0.6000 ;
    END
  END D[189]
  PIN D[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 325.8500 0.0000 325.9500 0.6000 ;
    END
  END D[188]
  PIN D[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 324.2500 0.0000 324.3500 0.6000 ;
    END
  END D[187]
  PIN D[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 322.6500 0.0000 322.7500 0.6000 ;
    END
  END D[186]
  PIN D[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 321.0500 0.0000 321.1500 0.6000 ;
    END
  END D[185]
  PIN D[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 319.4500 0.0000 319.5500 0.6000 ;
    END
  END D[184]
  PIN D[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 317.8500 0.0000 317.9500 0.6000 ;
    END
  END D[183]
  PIN D[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 316.2500 0.0000 316.3500 0.6000 ;
    END
  END D[182]
  PIN D[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 314.6500 0.0000 314.7500 0.6000 ;
    END
  END D[181]
  PIN D[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 313.0500 0.0000 313.1500 0.6000 ;
    END
  END D[180]
  PIN D[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 311.4500 0.0000 311.5500 0.6000 ;
    END
  END D[179]
  PIN D[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 309.8500 0.0000 309.9500 0.6000 ;
    END
  END D[178]
  PIN D[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 308.2500 0.0000 308.3500 0.6000 ;
    END
  END D[177]
  PIN D[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 306.6500 0.0000 306.7500 0.6000 ;
    END
  END D[176]
  PIN D[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 305.0500 0.0000 305.1500 0.6000 ;
    END
  END D[175]
  PIN D[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 303.4500 0.0000 303.5500 0.6000 ;
    END
  END D[174]
  PIN D[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 301.8500 0.0000 301.9500 0.6000 ;
    END
  END D[173]
  PIN D[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300.2500 0.0000 300.3500 0.6000 ;
    END
  END D[172]
  PIN D[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 298.6500 0.0000 298.7500 0.6000 ;
    END
  END D[171]
  PIN D[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 297.0500 0.0000 297.1500 0.6000 ;
    END
  END D[170]
  PIN D[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.4500 0.0000 295.5500 0.6000 ;
    END
  END D[169]
  PIN D[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 293.8500 0.0000 293.9500 0.6000 ;
    END
  END D[168]
  PIN D[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 292.2500 0.0000 292.3500 0.6000 ;
    END
  END D[167]
  PIN D[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 290.6500 0.0000 290.7500 0.6000 ;
    END
  END D[166]
  PIN D[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 289.0500 0.0000 289.1500 0.6000 ;
    END
  END D[165]
  PIN D[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 287.4500 0.0000 287.5500 0.6000 ;
    END
  END D[164]
  PIN D[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 285.8500 0.0000 285.9500 0.6000 ;
    END
  END D[163]
  PIN D[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 284.2500 0.0000 284.3500 0.6000 ;
    END
  END D[162]
  PIN D[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 282.6500 0.0000 282.7500 0.6000 ;
    END
  END D[161]
  PIN D[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 281.0500 0.0000 281.1500 0.6000 ;
    END
  END D[160]
  PIN D[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 279.4500 0.0000 279.5500 0.6000 ;
    END
  END D[159]
  PIN D[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 277.8500 0.0000 277.9500 0.6000 ;
    END
  END D[158]
  PIN D[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 276.2500 0.0000 276.3500 0.6000 ;
    END
  END D[157]
  PIN D[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 274.6500 0.0000 274.7500 0.6000 ;
    END
  END D[156]
  PIN D[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 273.0500 0.0000 273.1500 0.6000 ;
    END
  END D[155]
  PIN D[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 271.4500 0.0000 271.5500 0.6000 ;
    END
  END D[154]
  PIN D[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 269.8500 0.0000 269.9500 0.6000 ;
    END
  END D[153]
  PIN D[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 268.2500 0.0000 268.3500 0.6000 ;
    END
  END D[152]
  PIN D[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 266.6500 0.0000 266.7500 0.6000 ;
    END
  END D[151]
  PIN D[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 265.0500 0.0000 265.1500 0.6000 ;
    END
  END D[150]
  PIN D[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 263.4500 0.0000 263.5500 0.6000 ;
    END
  END D[149]
  PIN D[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 261.8500 0.0000 261.9500 0.6000 ;
    END
  END D[148]
  PIN D[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 260.2500 0.0000 260.3500 0.6000 ;
    END
  END D[147]
  PIN D[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 258.6500 0.0000 258.7500 0.6000 ;
    END
  END D[146]
  PIN D[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 257.0500 0.0000 257.1500 0.6000 ;
    END
  END D[145]
  PIN D[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 255.4500 0.0000 255.5500 0.6000 ;
    END
  END D[144]
  PIN D[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 253.8500 0.0000 253.9500 0.6000 ;
    END
  END D[143]
  PIN D[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 252.2500 0.0000 252.3500 0.6000 ;
    END
  END D[142]
  PIN D[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 250.6500 0.0000 250.7500 0.6000 ;
    END
  END D[141]
  PIN D[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 249.0500 0.0000 249.1500 0.6000 ;
    END
  END D[140]
  PIN D[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 247.4500 0.0000 247.5500 0.6000 ;
    END
  END D[139]
  PIN D[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 245.8500 0.0000 245.9500 0.6000 ;
    END
  END D[138]
  PIN D[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 244.2500 0.0000 244.3500 0.6000 ;
    END
  END D[137]
  PIN D[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 242.6500 0.0000 242.7500 0.6000 ;
    END
  END D[136]
  PIN D[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 241.0500 0.0000 241.1500 0.6000 ;
    END
  END D[135]
  PIN D[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 239.4500 0.0000 239.5500 0.6000 ;
    END
  END D[134]
  PIN D[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 237.8500 0.0000 237.9500 0.6000 ;
    END
  END D[133]
  PIN D[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 236.2500 0.0000 236.3500 0.6000 ;
    END
  END D[132]
  PIN D[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 234.6500 0.0000 234.7500 0.6000 ;
    END
  END D[131]
  PIN D[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 233.0500 0.0000 233.1500 0.6000 ;
    END
  END D[130]
  PIN D[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 231.4500 0.0000 231.5500 0.6000 ;
    END
  END D[129]
  PIN D[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 229.8500 0.0000 229.9500 0.6000 ;
    END
  END D[128]
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 228.2500 0.0000 228.3500 0.6000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 226.6500 0.0000 226.7500 0.6000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 225.0500 0.0000 225.1500 0.6000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 223.4500 0.0000 223.5500 0.6000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 221.8500 0.0000 221.9500 0.6000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220.2500 0.0000 220.3500 0.6000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 218.6500 0.0000 218.7500 0.6000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 217.0500 0.0000 217.1500 0.6000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 215.4500 0.0000 215.5500 0.6000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 213.8500 0.0000 213.9500 0.6000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 212.2500 0.0000 212.3500 0.6000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 210.6500 0.0000 210.7500 0.6000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 209.0500 0.0000 209.1500 0.6000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 207.4500 0.0000 207.5500 0.6000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 205.8500 0.0000 205.9500 0.6000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 204.2500 0.0000 204.3500 0.6000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 202.6500 0.0000 202.7500 0.6000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 201.0500 0.0000 201.1500 0.6000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 199.4500 0.0000 199.5500 0.6000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 197.8500 0.0000 197.9500 0.6000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 196.2500 0.0000 196.3500 0.6000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 194.6500 0.0000 194.7500 0.6000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 193.0500 0.0000 193.1500 0.6000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 191.4500 0.0000 191.5500 0.6000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 189.8500 0.0000 189.9500 0.6000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 188.2500 0.0000 188.3500 0.6000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 186.6500 0.0000 186.7500 0.6000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 185.0500 0.0000 185.1500 0.6000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.4500 0.0000 183.5500 0.6000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 181.8500 0.0000 181.9500 0.6000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.2500 0.0000 180.3500 0.6000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.6500 0.0000 178.7500 0.6000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.0500 0.0000 177.1500 0.6000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.4500 0.0000 175.5500 0.6000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.8500 0.0000 173.9500 0.6000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.2500 0.0000 172.3500 0.6000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 170.6500 0.0000 170.7500 0.6000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 169.0500 0.0000 169.1500 0.6000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.4500 0.0000 167.5500 0.6000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.8500 0.0000 165.9500 0.6000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.2500 0.0000 164.3500 0.6000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.6500 0.0000 162.7500 0.6000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.0500 0.0000 161.1500 0.6000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.4500 0.0000 159.5500 0.6000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 157.8500 0.0000 157.9500 0.6000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.2500 0.0000 156.3500 0.6000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.6500 0.0000 154.7500 0.6000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.0500 0.0000 153.1500 0.6000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.4500 0.0000 151.5500 0.6000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 149.8500 0.0000 149.9500 0.6000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.2500 0.0000 148.3500 0.6000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 146.6500 0.0000 146.7500 0.6000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 145.0500 0.0000 145.1500 0.6000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.4500 0.0000 143.5500 0.6000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.8500 0.0000 141.9500 0.6000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.2500 0.0000 140.3500 0.6000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.6500 0.0000 138.7500 0.6000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 137.0500 0.0000 137.1500 0.6000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.4500 0.0000 135.5500 0.6000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 133.8500 0.0000 133.9500 0.6000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.2500 0.0000 132.3500 0.6000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 130.6500 0.0000 130.7500 0.6000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.0500 0.0000 129.1500 0.6000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 127.4500 0.0000 127.5500 0.6000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.8500 0.0000 125.9500 0.6000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.2500 0.0000 124.3500 0.6000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.6500 0.0000 122.7500 0.6000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.0500 0.0000 121.1500 0.6000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.4500 0.0000 119.5500 0.6000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.8500 0.0000 117.9500 0.6000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.2500 0.0000 116.3500 0.6000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.6500 0.0000 114.7500 0.6000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.0500 0.0000 113.1500 0.6000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.4500 0.0000 111.5500 0.6000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.8500 0.0000 109.9500 0.6000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.2500 0.0000 108.3500 0.6000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.6500 0.0000 106.7500 0.6000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.0500 0.0000 105.1500 0.6000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.4500 0.0000 103.5500 0.6000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.8500 0.0000 101.9500 0.6000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.2500 0.0000 100.3500 0.6000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.6500 0.0000 98.7500 0.6000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.0500 0.0000 97.1500 0.6000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.4500 0.0000 95.5500 0.6000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.8500 0.0000 93.9500 0.6000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.2500 0.0000 92.3500 0.6000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.6500 0.0000 90.7500 0.6000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.0500 0.0000 89.1500 0.6000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.4500 0.0000 87.5500 0.6000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.8500 0.0000 85.9500 0.6000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.2500 0.0000 84.3500 0.6000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.6500 0.0000 82.7500 0.6000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.0500 0.0000 81.1500 0.6000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.4500 0.0000 79.5500 0.6000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 77.8500 0.0000 77.9500 0.6000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.2500 0.0000 76.3500 0.6000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 74.6500 0.0000 74.7500 0.6000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.0500 0.0000 73.1500 0.6000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.4500 0.0000 71.5500 0.6000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 69.8500 0.0000 69.9500 0.6000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.2500 0.0000 68.3500 0.6000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 66.6500 0.0000 66.7500 0.6000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.0500 0.0000 65.1500 0.6000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 63.4500 0.0000 63.5500 0.6000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 61.8500 0.0000 61.9500 0.6000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60.2500 0.0000 60.3500 0.6000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.6500 0.0000 58.7500 0.6000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 57.0500 0.0000 57.1500 0.6000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.4500 0.0000 55.5500 0.6000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 53.8500 0.0000 53.9500 0.6000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.2500 0.0000 52.3500 0.6000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 50.6500 0.0000 50.7500 0.6000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 49.0500 0.0000 49.1500 0.6000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 47.4500 0.0000 47.5500 0.6000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 45.8500 0.0000 45.9500 0.6000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 44.2500 0.0000 44.3500 0.6000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 42.6500 0.0000 42.7500 0.6000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 41.0500 0.0000 41.1500 0.6000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.4500 0.0000 39.5500 0.6000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 37.8500 0.0000 37.9500 0.6000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 36.2500 0.0000 36.3500 0.6000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 34.6500 0.0000 34.7500 0.6000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 33.0500 0.0000 33.1500 0.6000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 31.4500 0.0000 31.5500 0.6000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 29.8500 0.0000 29.9500 0.6000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 28.2500 0.0000 28.3500 0.6000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 26.6500 0.0000 26.7500 0.6000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 25.0500 0.0000 25.1500 0.6000 ;
    END
  END D[0]
  PIN Q[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 433.0500 102.2000 433.1500 102.8000 ;
    END
  END Q[255]
  PIN Q[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 431.4500 102.2000 431.5500 102.8000 ;
    END
  END Q[254]
  PIN Q[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 429.8500 102.2000 429.9500 102.8000 ;
    END
  END Q[253]
  PIN Q[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 428.2500 102.2000 428.3500 102.8000 ;
    END
  END Q[252]
  PIN Q[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 426.6500 102.2000 426.7500 102.8000 ;
    END
  END Q[251]
  PIN Q[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 425.0500 102.2000 425.1500 102.8000 ;
    END
  END Q[250]
  PIN Q[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 423.4500 102.2000 423.5500 102.8000 ;
    END
  END Q[249]
  PIN Q[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 421.8500 102.2000 421.9500 102.8000 ;
    END
  END Q[248]
  PIN Q[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 420.2500 102.2000 420.3500 102.8000 ;
    END
  END Q[247]
  PIN Q[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 418.6500 102.2000 418.7500 102.8000 ;
    END
  END Q[246]
  PIN Q[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 417.0500 102.2000 417.1500 102.8000 ;
    END
  END Q[245]
  PIN Q[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 415.4500 102.2000 415.5500 102.8000 ;
    END
  END Q[244]
  PIN Q[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 413.8500 102.2000 413.9500 102.8000 ;
    END
  END Q[243]
  PIN Q[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 412.2500 102.2000 412.3500 102.8000 ;
    END
  END Q[242]
  PIN Q[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 410.6500 102.2000 410.7500 102.8000 ;
    END
  END Q[241]
  PIN Q[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 409.0500 102.2000 409.1500 102.8000 ;
    END
  END Q[240]
  PIN Q[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 407.4500 102.2000 407.5500 102.8000 ;
    END
  END Q[239]
  PIN Q[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 405.8500 102.2000 405.9500 102.8000 ;
    END
  END Q[238]
  PIN Q[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 404.2500 102.2000 404.3500 102.8000 ;
    END
  END Q[237]
  PIN Q[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 402.6500 102.2000 402.7500 102.8000 ;
    END
  END Q[236]
  PIN Q[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.0500 102.2000 401.1500 102.8000 ;
    END
  END Q[235]
  PIN Q[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 399.4500 102.2000 399.5500 102.8000 ;
    END
  END Q[234]
  PIN Q[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 397.8500 102.2000 397.9500 102.8000 ;
    END
  END Q[233]
  PIN Q[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 396.2500 102.2000 396.3500 102.8000 ;
    END
  END Q[232]
  PIN Q[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 394.6500 102.2000 394.7500 102.8000 ;
    END
  END Q[231]
  PIN Q[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 393.0500 102.2000 393.1500 102.8000 ;
    END
  END Q[230]
  PIN Q[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 391.4500 102.2000 391.5500 102.8000 ;
    END
  END Q[229]
  PIN Q[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 389.8500 102.2000 389.9500 102.8000 ;
    END
  END Q[228]
  PIN Q[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 388.2500 102.2000 388.3500 102.8000 ;
    END
  END Q[227]
  PIN Q[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 386.6500 102.2000 386.7500 102.8000 ;
    END
  END Q[226]
  PIN Q[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 385.0500 102.2000 385.1500 102.8000 ;
    END
  END Q[225]
  PIN Q[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 383.4500 102.2000 383.5500 102.8000 ;
    END
  END Q[224]
  PIN Q[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 381.8500 102.2000 381.9500 102.8000 ;
    END
  END Q[223]
  PIN Q[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380.2500 102.2000 380.3500 102.8000 ;
    END
  END Q[222]
  PIN Q[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 378.6500 102.2000 378.7500 102.8000 ;
    END
  END Q[221]
  PIN Q[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 377.0500 102.2000 377.1500 102.8000 ;
    END
  END Q[220]
  PIN Q[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 375.4500 102.2000 375.5500 102.8000 ;
    END
  END Q[219]
  PIN Q[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 373.8500 102.2000 373.9500 102.8000 ;
    END
  END Q[218]
  PIN Q[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 372.2500 102.2000 372.3500 102.8000 ;
    END
  END Q[217]
  PIN Q[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 370.6500 102.2000 370.7500 102.8000 ;
    END
  END Q[216]
  PIN Q[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 369.0500 102.2000 369.1500 102.8000 ;
    END
  END Q[215]
  PIN Q[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 367.4500 102.2000 367.5500 102.8000 ;
    END
  END Q[214]
  PIN Q[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 365.8500 102.2000 365.9500 102.8000 ;
    END
  END Q[213]
  PIN Q[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 364.2500 102.2000 364.3500 102.8000 ;
    END
  END Q[212]
  PIN Q[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 362.6500 102.2000 362.7500 102.8000 ;
    END
  END Q[211]
  PIN Q[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 361.0500 102.2000 361.1500 102.8000 ;
    END
  END Q[210]
  PIN Q[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 359.4500 102.2000 359.5500 102.8000 ;
    END
  END Q[209]
  PIN Q[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 357.8500 102.2000 357.9500 102.8000 ;
    END
  END Q[208]
  PIN Q[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 356.2500 102.2000 356.3500 102.8000 ;
    END
  END Q[207]
  PIN Q[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 354.6500 102.2000 354.7500 102.8000 ;
    END
  END Q[206]
  PIN Q[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 353.0500 102.2000 353.1500 102.8000 ;
    END
  END Q[205]
  PIN Q[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 351.4500 102.2000 351.5500 102.8000 ;
    END
  END Q[204]
  PIN Q[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 349.8500 102.2000 349.9500 102.8000 ;
    END
  END Q[203]
  PIN Q[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 348.2500 102.2000 348.3500 102.8000 ;
    END
  END Q[202]
  PIN Q[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 346.6500 102.2000 346.7500 102.8000 ;
    END
  END Q[201]
  PIN Q[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 345.0500 102.2000 345.1500 102.8000 ;
    END
  END Q[200]
  PIN Q[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 343.4500 102.2000 343.5500 102.8000 ;
    END
  END Q[199]
  PIN Q[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 341.8500 102.2000 341.9500 102.8000 ;
    END
  END Q[198]
  PIN Q[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 340.2500 102.2000 340.3500 102.8000 ;
    END
  END Q[197]
  PIN Q[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 338.6500 102.2000 338.7500 102.8000 ;
    END
  END Q[196]
  PIN Q[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 337.0500 102.2000 337.1500 102.8000 ;
    END
  END Q[195]
  PIN Q[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 335.4500 102.2000 335.5500 102.8000 ;
    END
  END Q[194]
  PIN Q[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 333.8500 102.2000 333.9500 102.8000 ;
    END
  END Q[193]
  PIN Q[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 332.2500 102.2000 332.3500 102.8000 ;
    END
  END Q[192]
  PIN Q[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 330.6500 102.2000 330.7500 102.8000 ;
    END
  END Q[191]
  PIN Q[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 329.0500 102.2000 329.1500 102.8000 ;
    END
  END Q[190]
  PIN Q[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.4500 102.2000 327.5500 102.8000 ;
    END
  END Q[189]
  PIN Q[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 325.8500 102.2000 325.9500 102.8000 ;
    END
  END Q[188]
  PIN Q[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 324.2500 102.2000 324.3500 102.8000 ;
    END
  END Q[187]
  PIN Q[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 322.6500 102.2000 322.7500 102.8000 ;
    END
  END Q[186]
  PIN Q[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 321.0500 102.2000 321.1500 102.8000 ;
    END
  END Q[185]
  PIN Q[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 319.4500 102.2000 319.5500 102.8000 ;
    END
  END Q[184]
  PIN Q[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 317.8500 102.2000 317.9500 102.8000 ;
    END
  END Q[183]
  PIN Q[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 316.2500 102.2000 316.3500 102.8000 ;
    END
  END Q[182]
  PIN Q[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 314.6500 102.2000 314.7500 102.8000 ;
    END
  END Q[181]
  PIN Q[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 313.0500 102.2000 313.1500 102.8000 ;
    END
  END Q[180]
  PIN Q[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 311.4500 102.2000 311.5500 102.8000 ;
    END
  END Q[179]
  PIN Q[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 309.8500 102.2000 309.9500 102.8000 ;
    END
  END Q[178]
  PIN Q[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 308.2500 102.2000 308.3500 102.8000 ;
    END
  END Q[177]
  PIN Q[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 306.6500 102.2000 306.7500 102.8000 ;
    END
  END Q[176]
  PIN Q[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 305.0500 102.2000 305.1500 102.8000 ;
    END
  END Q[175]
  PIN Q[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 303.4500 102.2000 303.5500 102.8000 ;
    END
  END Q[174]
  PIN Q[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 301.8500 102.2000 301.9500 102.8000 ;
    END
  END Q[173]
  PIN Q[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300.2500 102.2000 300.3500 102.8000 ;
    END
  END Q[172]
  PIN Q[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 298.6500 102.2000 298.7500 102.8000 ;
    END
  END Q[171]
  PIN Q[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 297.0500 102.2000 297.1500 102.8000 ;
    END
  END Q[170]
  PIN Q[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.4500 102.2000 295.5500 102.8000 ;
    END
  END Q[169]
  PIN Q[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 293.8500 102.2000 293.9500 102.8000 ;
    END
  END Q[168]
  PIN Q[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 292.2500 102.2000 292.3500 102.8000 ;
    END
  END Q[167]
  PIN Q[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 290.6500 102.2000 290.7500 102.8000 ;
    END
  END Q[166]
  PIN Q[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 289.0500 102.2000 289.1500 102.8000 ;
    END
  END Q[165]
  PIN Q[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 287.4500 102.2000 287.5500 102.8000 ;
    END
  END Q[164]
  PIN Q[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 285.8500 102.2000 285.9500 102.8000 ;
    END
  END Q[163]
  PIN Q[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 284.2500 102.2000 284.3500 102.8000 ;
    END
  END Q[162]
  PIN Q[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 282.6500 102.2000 282.7500 102.8000 ;
    END
  END Q[161]
  PIN Q[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 281.0500 102.2000 281.1500 102.8000 ;
    END
  END Q[160]
  PIN Q[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 279.4500 102.2000 279.5500 102.8000 ;
    END
  END Q[159]
  PIN Q[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 277.8500 102.2000 277.9500 102.8000 ;
    END
  END Q[158]
  PIN Q[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 276.2500 102.2000 276.3500 102.8000 ;
    END
  END Q[157]
  PIN Q[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 274.6500 102.2000 274.7500 102.8000 ;
    END
  END Q[156]
  PIN Q[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 273.0500 102.2000 273.1500 102.8000 ;
    END
  END Q[155]
  PIN Q[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 271.4500 102.2000 271.5500 102.8000 ;
    END
  END Q[154]
  PIN Q[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 269.8500 102.2000 269.9500 102.8000 ;
    END
  END Q[153]
  PIN Q[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 268.2500 102.2000 268.3500 102.8000 ;
    END
  END Q[152]
  PIN Q[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 266.6500 102.2000 266.7500 102.8000 ;
    END
  END Q[151]
  PIN Q[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 265.0500 102.2000 265.1500 102.8000 ;
    END
  END Q[150]
  PIN Q[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 263.4500 102.2000 263.5500 102.8000 ;
    END
  END Q[149]
  PIN Q[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 261.8500 102.2000 261.9500 102.8000 ;
    END
  END Q[148]
  PIN Q[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 260.2500 102.2000 260.3500 102.8000 ;
    END
  END Q[147]
  PIN Q[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 258.6500 102.2000 258.7500 102.8000 ;
    END
  END Q[146]
  PIN Q[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 257.0500 102.2000 257.1500 102.8000 ;
    END
  END Q[145]
  PIN Q[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 255.4500 102.2000 255.5500 102.8000 ;
    END
  END Q[144]
  PIN Q[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 253.8500 102.2000 253.9500 102.8000 ;
    END
  END Q[143]
  PIN Q[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 252.2500 102.2000 252.3500 102.8000 ;
    END
  END Q[142]
  PIN Q[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 250.6500 102.2000 250.7500 102.8000 ;
    END
  END Q[141]
  PIN Q[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 249.0500 102.2000 249.1500 102.8000 ;
    END
  END Q[140]
  PIN Q[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 247.4500 102.2000 247.5500 102.8000 ;
    END
  END Q[139]
  PIN Q[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 245.8500 102.2000 245.9500 102.8000 ;
    END
  END Q[138]
  PIN Q[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 244.2500 102.2000 244.3500 102.8000 ;
    END
  END Q[137]
  PIN Q[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 242.6500 102.2000 242.7500 102.8000 ;
    END
  END Q[136]
  PIN Q[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 241.0500 102.2000 241.1500 102.8000 ;
    END
  END Q[135]
  PIN Q[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 239.4500 102.2000 239.5500 102.8000 ;
    END
  END Q[134]
  PIN Q[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 237.8500 102.2000 237.9500 102.8000 ;
    END
  END Q[133]
  PIN Q[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 236.2500 102.2000 236.3500 102.8000 ;
    END
  END Q[132]
  PIN Q[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 234.6500 102.2000 234.7500 102.8000 ;
    END
  END Q[131]
  PIN Q[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 233.0500 102.2000 233.1500 102.8000 ;
    END
  END Q[130]
  PIN Q[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 231.4500 102.2000 231.5500 102.8000 ;
    END
  END Q[129]
  PIN Q[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 229.8500 102.2000 229.9500 102.8000 ;
    END
  END Q[128]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 228.2500 102.2000 228.3500 102.8000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 226.6500 102.2000 226.7500 102.8000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 225.0500 102.2000 225.1500 102.8000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 223.4500 102.2000 223.5500 102.8000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 221.8500 102.2000 221.9500 102.8000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220.2500 102.2000 220.3500 102.8000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 218.6500 102.2000 218.7500 102.8000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 217.0500 102.2000 217.1500 102.8000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 215.4500 102.2000 215.5500 102.8000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 213.8500 102.2000 213.9500 102.8000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 212.2500 102.2000 212.3500 102.8000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 210.6500 102.2000 210.7500 102.8000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 209.0500 102.2000 209.1500 102.8000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 207.4500 102.2000 207.5500 102.8000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 205.8500 102.2000 205.9500 102.8000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 204.2500 102.2000 204.3500 102.8000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 202.6500 102.2000 202.7500 102.8000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 201.0500 102.2000 201.1500 102.8000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 199.4500 102.2000 199.5500 102.8000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 197.8500 102.2000 197.9500 102.8000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 196.2500 102.2000 196.3500 102.8000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 194.6500 102.2000 194.7500 102.8000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 193.0500 102.2000 193.1500 102.8000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 191.4500 102.2000 191.5500 102.8000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 189.8500 102.2000 189.9500 102.8000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 188.2500 102.2000 188.3500 102.8000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 186.6500 102.2000 186.7500 102.8000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 185.0500 102.2000 185.1500 102.8000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.4500 102.2000 183.5500 102.8000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 181.8500 102.2000 181.9500 102.8000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.2500 102.2000 180.3500 102.8000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.6500 102.2000 178.7500 102.8000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.0500 102.2000 177.1500 102.8000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.4500 102.2000 175.5500 102.8000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.8500 102.2000 173.9500 102.8000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.2500 102.2000 172.3500 102.8000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 170.6500 102.2000 170.7500 102.8000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 169.0500 102.2000 169.1500 102.8000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.4500 102.2000 167.5500 102.8000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.8500 102.2000 165.9500 102.8000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.2500 102.2000 164.3500 102.8000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.6500 102.2000 162.7500 102.8000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.0500 102.2000 161.1500 102.8000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.4500 102.2000 159.5500 102.8000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 157.8500 102.2000 157.9500 102.8000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.2500 102.2000 156.3500 102.8000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.6500 102.2000 154.7500 102.8000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.0500 102.2000 153.1500 102.8000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.4500 102.2000 151.5500 102.8000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 149.8500 102.2000 149.9500 102.8000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.2500 102.2000 148.3500 102.8000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 146.6500 102.2000 146.7500 102.8000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 145.0500 102.2000 145.1500 102.8000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.4500 102.2000 143.5500 102.8000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.8500 102.2000 141.9500 102.8000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.2500 102.2000 140.3500 102.8000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.6500 102.2000 138.7500 102.8000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 137.0500 102.2000 137.1500 102.8000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.4500 102.2000 135.5500 102.8000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 133.8500 102.2000 133.9500 102.8000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.2500 102.2000 132.3500 102.8000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 130.6500 102.2000 130.7500 102.8000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.0500 102.2000 129.1500 102.8000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 127.4500 102.2000 127.5500 102.8000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.8500 102.2000 125.9500 102.8000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.2500 102.2000 124.3500 102.8000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.6500 102.2000 122.7500 102.8000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.0500 102.2000 121.1500 102.8000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.4500 102.2000 119.5500 102.8000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.8500 102.2000 117.9500 102.8000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.2500 102.2000 116.3500 102.8000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.6500 102.2000 114.7500 102.8000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.0500 102.2000 113.1500 102.8000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.4500 102.2000 111.5500 102.8000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.8500 102.2000 109.9500 102.8000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.2500 102.2000 108.3500 102.8000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.6500 102.2000 106.7500 102.8000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.0500 102.2000 105.1500 102.8000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.4500 102.2000 103.5500 102.8000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.8500 102.2000 101.9500 102.8000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.2500 102.2000 100.3500 102.8000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.6500 102.2000 98.7500 102.8000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.0500 102.2000 97.1500 102.8000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.4500 102.2000 95.5500 102.8000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.8500 102.2000 93.9500 102.8000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.2500 102.2000 92.3500 102.8000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.6500 102.2000 90.7500 102.8000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.0500 102.2000 89.1500 102.8000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.4500 102.2000 87.5500 102.8000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.8500 102.2000 85.9500 102.8000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.2500 102.2000 84.3500 102.8000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.6500 102.2000 82.7500 102.8000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.0500 102.2000 81.1500 102.8000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.4500 102.2000 79.5500 102.8000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 77.8500 102.2000 77.9500 102.8000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.2500 102.2000 76.3500 102.8000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 74.6500 102.2000 74.7500 102.8000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.0500 102.2000 73.1500 102.8000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.4500 102.2000 71.5500 102.8000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 69.8500 102.2000 69.9500 102.8000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.2500 102.2000 68.3500 102.8000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 66.6500 102.2000 66.7500 102.8000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.0500 102.2000 65.1500 102.8000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 63.4500 102.2000 63.5500 102.8000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 61.8500 102.2000 61.9500 102.8000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60.2500 102.2000 60.3500 102.8000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.6500 102.2000 58.7500 102.8000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 57.0500 102.2000 57.1500 102.8000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.4500 102.2000 55.5500 102.8000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 53.8500 102.2000 53.9500 102.8000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.2500 102.2000 52.3500 102.8000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 50.6500 102.2000 50.7500 102.8000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 49.0500 102.2000 49.1500 102.8000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 47.4500 102.2000 47.5500 102.8000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 45.8500 102.2000 45.9500 102.8000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 44.2500 102.2000 44.3500 102.8000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 42.6500 102.2000 42.7500 102.8000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 41.0500 102.2000 41.1500 102.8000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.4500 102.2000 39.5500 102.8000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 37.8500 102.2000 37.9500 102.8000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 36.2500 102.2000 36.3500 102.8000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 34.6500 102.2000 34.7500 102.8000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 33.0500 102.2000 33.1500 102.8000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 31.4500 102.2000 31.5500 102.8000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 29.8500 102.2000 29.9500 102.8000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 28.2500 102.2000 28.3500 102.8000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 26.6500 102.2000 26.7500 102.8000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 25.0500 102.2000 25.1500 102.8000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 47.5500 0.6000 47.6500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 39.5500 0.6000 39.6500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 51.5500 0.6000 51.6500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.5500 0.6000 55.6500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 59.5500 0.6000 59.6500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 63.5500 0.6000 63.6500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 157.0650 10.0000 159.0650 92.8000 ;
        RECT 30.0000 10.0000 32.0000 92.8000 ;
        RECT 411.1950 10.0000 413.1950 92.8000 ;
        RECT 284.1300 10.0000 286.1300 92.8000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 164.0650 10.0000 166.0650 92.8000 ;
        RECT 37.0000 10.0000 39.0000 92.8000 ;
        RECT 418.1950 10.0000 420.1950 92.8000 ;
        RECT 291.1300 10.0000 293.1300 92.8000 ;
        RECT 37.0000 9.8350 39.0000 10.1650 ;
        RECT 164.0650 9.8350 166.0650 10.1650 ;
        RECT 291.1300 9.8350 293.1300 10.1650 ;
        RECT 418.1950 9.8350 420.1950 10.1650 ;
        RECT 37.0000 92.6350 39.0000 92.9650 ;
        RECT 164.0650 92.6350 166.0650 92.9650 ;
        RECT 291.1300 92.6350 293.1300 92.9650 ;
        RECT 418.1950 92.6350 420.1950 92.9650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 450.2000 102.8000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 450.2000 102.8000 ;
    LAYER M3 ;
      RECT 433.3100 102.0400 450.2000 102.8000 ;
      RECT 431.7100 102.0400 432.8900 102.8000 ;
      RECT 430.1100 102.0400 431.2900 102.8000 ;
      RECT 428.5100 102.0400 429.6900 102.8000 ;
      RECT 426.9100 102.0400 428.0900 102.8000 ;
      RECT 425.3100 102.0400 426.4900 102.8000 ;
      RECT 423.7100 102.0400 424.8900 102.8000 ;
      RECT 422.1100 102.0400 423.2900 102.8000 ;
      RECT 420.5100 102.0400 421.6900 102.8000 ;
      RECT 418.9100 102.0400 420.0900 102.8000 ;
      RECT 417.3100 102.0400 418.4900 102.8000 ;
      RECT 415.7100 102.0400 416.8900 102.8000 ;
      RECT 414.1100 102.0400 415.2900 102.8000 ;
      RECT 412.5100 102.0400 413.6900 102.8000 ;
      RECT 410.9100 102.0400 412.0900 102.8000 ;
      RECT 409.3100 102.0400 410.4900 102.8000 ;
      RECT 407.7100 102.0400 408.8900 102.8000 ;
      RECT 406.1100 102.0400 407.2900 102.8000 ;
      RECT 404.5100 102.0400 405.6900 102.8000 ;
      RECT 402.9100 102.0400 404.0900 102.8000 ;
      RECT 401.3100 102.0400 402.4900 102.8000 ;
      RECT 399.7100 102.0400 400.8900 102.8000 ;
      RECT 398.1100 102.0400 399.2900 102.8000 ;
      RECT 396.5100 102.0400 397.6900 102.8000 ;
      RECT 394.9100 102.0400 396.0900 102.8000 ;
      RECT 393.3100 102.0400 394.4900 102.8000 ;
      RECT 391.7100 102.0400 392.8900 102.8000 ;
      RECT 390.1100 102.0400 391.2900 102.8000 ;
      RECT 388.5100 102.0400 389.6900 102.8000 ;
      RECT 386.9100 102.0400 388.0900 102.8000 ;
      RECT 385.3100 102.0400 386.4900 102.8000 ;
      RECT 383.7100 102.0400 384.8900 102.8000 ;
      RECT 382.1100 102.0400 383.2900 102.8000 ;
      RECT 380.5100 102.0400 381.6900 102.8000 ;
      RECT 378.9100 102.0400 380.0900 102.8000 ;
      RECT 377.3100 102.0400 378.4900 102.8000 ;
      RECT 375.7100 102.0400 376.8900 102.8000 ;
      RECT 374.1100 102.0400 375.2900 102.8000 ;
      RECT 372.5100 102.0400 373.6900 102.8000 ;
      RECT 370.9100 102.0400 372.0900 102.8000 ;
      RECT 369.3100 102.0400 370.4900 102.8000 ;
      RECT 367.7100 102.0400 368.8900 102.8000 ;
      RECT 366.1100 102.0400 367.2900 102.8000 ;
      RECT 364.5100 102.0400 365.6900 102.8000 ;
      RECT 362.9100 102.0400 364.0900 102.8000 ;
      RECT 361.3100 102.0400 362.4900 102.8000 ;
      RECT 359.7100 102.0400 360.8900 102.8000 ;
      RECT 358.1100 102.0400 359.2900 102.8000 ;
      RECT 356.5100 102.0400 357.6900 102.8000 ;
      RECT 354.9100 102.0400 356.0900 102.8000 ;
      RECT 353.3100 102.0400 354.4900 102.8000 ;
      RECT 351.7100 102.0400 352.8900 102.8000 ;
      RECT 350.1100 102.0400 351.2900 102.8000 ;
      RECT 348.5100 102.0400 349.6900 102.8000 ;
      RECT 346.9100 102.0400 348.0900 102.8000 ;
      RECT 345.3100 102.0400 346.4900 102.8000 ;
      RECT 343.7100 102.0400 344.8900 102.8000 ;
      RECT 342.1100 102.0400 343.2900 102.8000 ;
      RECT 340.5100 102.0400 341.6900 102.8000 ;
      RECT 338.9100 102.0400 340.0900 102.8000 ;
      RECT 337.3100 102.0400 338.4900 102.8000 ;
      RECT 335.7100 102.0400 336.8900 102.8000 ;
      RECT 334.1100 102.0400 335.2900 102.8000 ;
      RECT 332.5100 102.0400 333.6900 102.8000 ;
      RECT 330.9100 102.0400 332.0900 102.8000 ;
      RECT 329.3100 102.0400 330.4900 102.8000 ;
      RECT 327.7100 102.0400 328.8900 102.8000 ;
      RECT 326.1100 102.0400 327.2900 102.8000 ;
      RECT 324.5100 102.0400 325.6900 102.8000 ;
      RECT 322.9100 102.0400 324.0900 102.8000 ;
      RECT 321.3100 102.0400 322.4900 102.8000 ;
      RECT 319.7100 102.0400 320.8900 102.8000 ;
      RECT 318.1100 102.0400 319.2900 102.8000 ;
      RECT 316.5100 102.0400 317.6900 102.8000 ;
      RECT 314.9100 102.0400 316.0900 102.8000 ;
      RECT 313.3100 102.0400 314.4900 102.8000 ;
      RECT 311.7100 102.0400 312.8900 102.8000 ;
      RECT 310.1100 102.0400 311.2900 102.8000 ;
      RECT 308.5100 102.0400 309.6900 102.8000 ;
      RECT 306.9100 102.0400 308.0900 102.8000 ;
      RECT 305.3100 102.0400 306.4900 102.8000 ;
      RECT 303.7100 102.0400 304.8900 102.8000 ;
      RECT 302.1100 102.0400 303.2900 102.8000 ;
      RECT 300.5100 102.0400 301.6900 102.8000 ;
      RECT 298.9100 102.0400 300.0900 102.8000 ;
      RECT 297.3100 102.0400 298.4900 102.8000 ;
      RECT 295.7100 102.0400 296.8900 102.8000 ;
      RECT 294.1100 102.0400 295.2900 102.8000 ;
      RECT 292.5100 102.0400 293.6900 102.8000 ;
      RECT 290.9100 102.0400 292.0900 102.8000 ;
      RECT 289.3100 102.0400 290.4900 102.8000 ;
      RECT 287.7100 102.0400 288.8900 102.8000 ;
      RECT 286.1100 102.0400 287.2900 102.8000 ;
      RECT 284.5100 102.0400 285.6900 102.8000 ;
      RECT 282.9100 102.0400 284.0900 102.8000 ;
      RECT 281.3100 102.0400 282.4900 102.8000 ;
      RECT 279.7100 102.0400 280.8900 102.8000 ;
      RECT 278.1100 102.0400 279.2900 102.8000 ;
      RECT 276.5100 102.0400 277.6900 102.8000 ;
      RECT 274.9100 102.0400 276.0900 102.8000 ;
      RECT 273.3100 102.0400 274.4900 102.8000 ;
      RECT 271.7100 102.0400 272.8900 102.8000 ;
      RECT 270.1100 102.0400 271.2900 102.8000 ;
      RECT 268.5100 102.0400 269.6900 102.8000 ;
      RECT 266.9100 102.0400 268.0900 102.8000 ;
      RECT 265.3100 102.0400 266.4900 102.8000 ;
      RECT 263.7100 102.0400 264.8900 102.8000 ;
      RECT 262.1100 102.0400 263.2900 102.8000 ;
      RECT 260.5100 102.0400 261.6900 102.8000 ;
      RECT 258.9100 102.0400 260.0900 102.8000 ;
      RECT 257.3100 102.0400 258.4900 102.8000 ;
      RECT 255.7100 102.0400 256.8900 102.8000 ;
      RECT 254.1100 102.0400 255.2900 102.8000 ;
      RECT 252.5100 102.0400 253.6900 102.8000 ;
      RECT 250.9100 102.0400 252.0900 102.8000 ;
      RECT 249.3100 102.0400 250.4900 102.8000 ;
      RECT 247.7100 102.0400 248.8900 102.8000 ;
      RECT 246.1100 102.0400 247.2900 102.8000 ;
      RECT 244.5100 102.0400 245.6900 102.8000 ;
      RECT 242.9100 102.0400 244.0900 102.8000 ;
      RECT 241.3100 102.0400 242.4900 102.8000 ;
      RECT 239.7100 102.0400 240.8900 102.8000 ;
      RECT 238.1100 102.0400 239.2900 102.8000 ;
      RECT 236.5100 102.0400 237.6900 102.8000 ;
      RECT 234.9100 102.0400 236.0900 102.8000 ;
      RECT 233.3100 102.0400 234.4900 102.8000 ;
      RECT 231.7100 102.0400 232.8900 102.8000 ;
      RECT 230.1100 102.0400 231.2900 102.8000 ;
      RECT 228.5100 102.0400 229.6900 102.8000 ;
      RECT 226.9100 102.0400 228.0900 102.8000 ;
      RECT 225.3100 102.0400 226.4900 102.8000 ;
      RECT 223.7100 102.0400 224.8900 102.8000 ;
      RECT 222.1100 102.0400 223.2900 102.8000 ;
      RECT 220.5100 102.0400 221.6900 102.8000 ;
      RECT 218.9100 102.0400 220.0900 102.8000 ;
      RECT 217.3100 102.0400 218.4900 102.8000 ;
      RECT 215.7100 102.0400 216.8900 102.8000 ;
      RECT 214.1100 102.0400 215.2900 102.8000 ;
      RECT 212.5100 102.0400 213.6900 102.8000 ;
      RECT 210.9100 102.0400 212.0900 102.8000 ;
      RECT 209.3100 102.0400 210.4900 102.8000 ;
      RECT 207.7100 102.0400 208.8900 102.8000 ;
      RECT 206.1100 102.0400 207.2900 102.8000 ;
      RECT 204.5100 102.0400 205.6900 102.8000 ;
      RECT 202.9100 102.0400 204.0900 102.8000 ;
      RECT 201.3100 102.0400 202.4900 102.8000 ;
      RECT 199.7100 102.0400 200.8900 102.8000 ;
      RECT 198.1100 102.0400 199.2900 102.8000 ;
      RECT 196.5100 102.0400 197.6900 102.8000 ;
      RECT 194.9100 102.0400 196.0900 102.8000 ;
      RECT 193.3100 102.0400 194.4900 102.8000 ;
      RECT 191.7100 102.0400 192.8900 102.8000 ;
      RECT 190.1100 102.0400 191.2900 102.8000 ;
      RECT 188.5100 102.0400 189.6900 102.8000 ;
      RECT 186.9100 102.0400 188.0900 102.8000 ;
      RECT 185.3100 102.0400 186.4900 102.8000 ;
      RECT 183.7100 102.0400 184.8900 102.8000 ;
      RECT 182.1100 102.0400 183.2900 102.8000 ;
      RECT 180.5100 102.0400 181.6900 102.8000 ;
      RECT 178.9100 102.0400 180.0900 102.8000 ;
      RECT 177.3100 102.0400 178.4900 102.8000 ;
      RECT 175.7100 102.0400 176.8900 102.8000 ;
      RECT 174.1100 102.0400 175.2900 102.8000 ;
      RECT 172.5100 102.0400 173.6900 102.8000 ;
      RECT 170.9100 102.0400 172.0900 102.8000 ;
      RECT 169.3100 102.0400 170.4900 102.8000 ;
      RECT 167.7100 102.0400 168.8900 102.8000 ;
      RECT 166.1100 102.0400 167.2900 102.8000 ;
      RECT 164.5100 102.0400 165.6900 102.8000 ;
      RECT 162.9100 102.0400 164.0900 102.8000 ;
      RECT 161.3100 102.0400 162.4900 102.8000 ;
      RECT 159.7100 102.0400 160.8900 102.8000 ;
      RECT 158.1100 102.0400 159.2900 102.8000 ;
      RECT 156.5100 102.0400 157.6900 102.8000 ;
      RECT 154.9100 102.0400 156.0900 102.8000 ;
      RECT 153.3100 102.0400 154.4900 102.8000 ;
      RECT 151.7100 102.0400 152.8900 102.8000 ;
      RECT 150.1100 102.0400 151.2900 102.8000 ;
      RECT 148.5100 102.0400 149.6900 102.8000 ;
      RECT 146.9100 102.0400 148.0900 102.8000 ;
      RECT 145.3100 102.0400 146.4900 102.8000 ;
      RECT 143.7100 102.0400 144.8900 102.8000 ;
      RECT 142.1100 102.0400 143.2900 102.8000 ;
      RECT 140.5100 102.0400 141.6900 102.8000 ;
      RECT 138.9100 102.0400 140.0900 102.8000 ;
      RECT 137.3100 102.0400 138.4900 102.8000 ;
      RECT 135.7100 102.0400 136.8900 102.8000 ;
      RECT 134.1100 102.0400 135.2900 102.8000 ;
      RECT 132.5100 102.0400 133.6900 102.8000 ;
      RECT 130.9100 102.0400 132.0900 102.8000 ;
      RECT 129.3100 102.0400 130.4900 102.8000 ;
      RECT 127.7100 102.0400 128.8900 102.8000 ;
      RECT 126.1100 102.0400 127.2900 102.8000 ;
      RECT 124.5100 102.0400 125.6900 102.8000 ;
      RECT 122.9100 102.0400 124.0900 102.8000 ;
      RECT 121.3100 102.0400 122.4900 102.8000 ;
      RECT 119.7100 102.0400 120.8900 102.8000 ;
      RECT 118.1100 102.0400 119.2900 102.8000 ;
      RECT 116.5100 102.0400 117.6900 102.8000 ;
      RECT 114.9100 102.0400 116.0900 102.8000 ;
      RECT 113.3100 102.0400 114.4900 102.8000 ;
      RECT 111.7100 102.0400 112.8900 102.8000 ;
      RECT 110.1100 102.0400 111.2900 102.8000 ;
      RECT 108.5100 102.0400 109.6900 102.8000 ;
      RECT 106.9100 102.0400 108.0900 102.8000 ;
      RECT 105.3100 102.0400 106.4900 102.8000 ;
      RECT 103.7100 102.0400 104.8900 102.8000 ;
      RECT 102.1100 102.0400 103.2900 102.8000 ;
      RECT 100.5100 102.0400 101.6900 102.8000 ;
      RECT 98.9100 102.0400 100.0900 102.8000 ;
      RECT 97.3100 102.0400 98.4900 102.8000 ;
      RECT 95.7100 102.0400 96.8900 102.8000 ;
      RECT 94.1100 102.0400 95.2900 102.8000 ;
      RECT 92.5100 102.0400 93.6900 102.8000 ;
      RECT 90.9100 102.0400 92.0900 102.8000 ;
      RECT 89.3100 102.0400 90.4900 102.8000 ;
      RECT 87.7100 102.0400 88.8900 102.8000 ;
      RECT 86.1100 102.0400 87.2900 102.8000 ;
      RECT 84.5100 102.0400 85.6900 102.8000 ;
      RECT 82.9100 102.0400 84.0900 102.8000 ;
      RECT 81.3100 102.0400 82.4900 102.8000 ;
      RECT 79.7100 102.0400 80.8900 102.8000 ;
      RECT 78.1100 102.0400 79.2900 102.8000 ;
      RECT 76.5100 102.0400 77.6900 102.8000 ;
      RECT 74.9100 102.0400 76.0900 102.8000 ;
      RECT 73.3100 102.0400 74.4900 102.8000 ;
      RECT 71.7100 102.0400 72.8900 102.8000 ;
      RECT 70.1100 102.0400 71.2900 102.8000 ;
      RECT 68.5100 102.0400 69.6900 102.8000 ;
      RECT 66.9100 102.0400 68.0900 102.8000 ;
      RECT 65.3100 102.0400 66.4900 102.8000 ;
      RECT 63.7100 102.0400 64.8900 102.8000 ;
      RECT 62.1100 102.0400 63.2900 102.8000 ;
      RECT 60.5100 102.0400 61.6900 102.8000 ;
      RECT 58.9100 102.0400 60.0900 102.8000 ;
      RECT 57.3100 102.0400 58.4900 102.8000 ;
      RECT 55.7100 102.0400 56.8900 102.8000 ;
      RECT 54.1100 102.0400 55.2900 102.8000 ;
      RECT 52.5100 102.0400 53.6900 102.8000 ;
      RECT 50.9100 102.0400 52.0900 102.8000 ;
      RECT 49.3100 102.0400 50.4900 102.8000 ;
      RECT 47.7100 102.0400 48.8900 102.8000 ;
      RECT 46.1100 102.0400 47.2900 102.8000 ;
      RECT 44.5100 102.0400 45.6900 102.8000 ;
      RECT 42.9100 102.0400 44.0900 102.8000 ;
      RECT 41.3100 102.0400 42.4900 102.8000 ;
      RECT 39.7100 102.0400 40.8900 102.8000 ;
      RECT 38.1100 102.0400 39.2900 102.8000 ;
      RECT 36.5100 102.0400 37.6900 102.8000 ;
      RECT 34.9100 102.0400 36.0900 102.8000 ;
      RECT 33.3100 102.0400 34.4900 102.8000 ;
      RECT 31.7100 102.0400 32.8900 102.8000 ;
      RECT 30.1100 102.0400 31.2900 102.8000 ;
      RECT 28.5100 102.0400 29.6900 102.8000 ;
      RECT 26.9100 102.0400 28.0900 102.8000 ;
      RECT 25.3100 102.0400 26.4900 102.8000 ;
      RECT 0.0000 102.0400 24.8900 102.8000 ;
      RECT 0.0000 63.7500 450.2000 102.0400 ;
      RECT 0.7000 63.4500 450.2000 63.7500 ;
      RECT 0.0000 59.7500 450.2000 63.4500 ;
      RECT 0.7000 59.4500 450.2000 59.7500 ;
      RECT 0.0000 55.7500 450.2000 59.4500 ;
      RECT 0.7000 55.4500 450.2000 55.7500 ;
      RECT 0.0000 51.7500 450.2000 55.4500 ;
      RECT 0.7000 51.4500 450.2000 51.7500 ;
      RECT 0.0000 47.7500 450.2000 51.4500 ;
      RECT 0.7000 47.4500 450.2000 47.7500 ;
      RECT 0.0000 43.7500 450.2000 47.4500 ;
      RECT 0.7000 43.4500 450.2000 43.7500 ;
      RECT 0.0000 39.7500 450.2000 43.4500 ;
      RECT 0.7000 39.4500 450.2000 39.7500 ;
      RECT 0.0000 0.7600 450.2000 39.4500 ;
      RECT 433.3100 0.0000 450.2000 0.7600 ;
      RECT 431.7100 0.0000 432.8900 0.7600 ;
      RECT 430.1100 0.0000 431.2900 0.7600 ;
      RECT 428.5100 0.0000 429.6900 0.7600 ;
      RECT 426.9100 0.0000 428.0900 0.7600 ;
      RECT 425.3100 0.0000 426.4900 0.7600 ;
      RECT 423.7100 0.0000 424.8900 0.7600 ;
      RECT 422.1100 0.0000 423.2900 0.7600 ;
      RECT 420.5100 0.0000 421.6900 0.7600 ;
      RECT 418.9100 0.0000 420.0900 0.7600 ;
      RECT 417.3100 0.0000 418.4900 0.7600 ;
      RECT 415.7100 0.0000 416.8900 0.7600 ;
      RECT 414.1100 0.0000 415.2900 0.7600 ;
      RECT 412.5100 0.0000 413.6900 0.7600 ;
      RECT 410.9100 0.0000 412.0900 0.7600 ;
      RECT 409.3100 0.0000 410.4900 0.7600 ;
      RECT 407.7100 0.0000 408.8900 0.7600 ;
      RECT 406.1100 0.0000 407.2900 0.7600 ;
      RECT 404.5100 0.0000 405.6900 0.7600 ;
      RECT 402.9100 0.0000 404.0900 0.7600 ;
      RECT 401.3100 0.0000 402.4900 0.7600 ;
      RECT 399.7100 0.0000 400.8900 0.7600 ;
      RECT 398.1100 0.0000 399.2900 0.7600 ;
      RECT 396.5100 0.0000 397.6900 0.7600 ;
      RECT 394.9100 0.0000 396.0900 0.7600 ;
      RECT 393.3100 0.0000 394.4900 0.7600 ;
      RECT 391.7100 0.0000 392.8900 0.7600 ;
      RECT 390.1100 0.0000 391.2900 0.7600 ;
      RECT 388.5100 0.0000 389.6900 0.7600 ;
      RECT 386.9100 0.0000 388.0900 0.7600 ;
      RECT 385.3100 0.0000 386.4900 0.7600 ;
      RECT 383.7100 0.0000 384.8900 0.7600 ;
      RECT 382.1100 0.0000 383.2900 0.7600 ;
      RECT 380.5100 0.0000 381.6900 0.7600 ;
      RECT 378.9100 0.0000 380.0900 0.7600 ;
      RECT 377.3100 0.0000 378.4900 0.7600 ;
      RECT 375.7100 0.0000 376.8900 0.7600 ;
      RECT 374.1100 0.0000 375.2900 0.7600 ;
      RECT 372.5100 0.0000 373.6900 0.7600 ;
      RECT 370.9100 0.0000 372.0900 0.7600 ;
      RECT 369.3100 0.0000 370.4900 0.7600 ;
      RECT 367.7100 0.0000 368.8900 0.7600 ;
      RECT 366.1100 0.0000 367.2900 0.7600 ;
      RECT 364.5100 0.0000 365.6900 0.7600 ;
      RECT 362.9100 0.0000 364.0900 0.7600 ;
      RECT 361.3100 0.0000 362.4900 0.7600 ;
      RECT 359.7100 0.0000 360.8900 0.7600 ;
      RECT 358.1100 0.0000 359.2900 0.7600 ;
      RECT 356.5100 0.0000 357.6900 0.7600 ;
      RECT 354.9100 0.0000 356.0900 0.7600 ;
      RECT 353.3100 0.0000 354.4900 0.7600 ;
      RECT 351.7100 0.0000 352.8900 0.7600 ;
      RECT 350.1100 0.0000 351.2900 0.7600 ;
      RECT 348.5100 0.0000 349.6900 0.7600 ;
      RECT 346.9100 0.0000 348.0900 0.7600 ;
      RECT 345.3100 0.0000 346.4900 0.7600 ;
      RECT 343.7100 0.0000 344.8900 0.7600 ;
      RECT 342.1100 0.0000 343.2900 0.7600 ;
      RECT 340.5100 0.0000 341.6900 0.7600 ;
      RECT 338.9100 0.0000 340.0900 0.7600 ;
      RECT 337.3100 0.0000 338.4900 0.7600 ;
      RECT 335.7100 0.0000 336.8900 0.7600 ;
      RECT 334.1100 0.0000 335.2900 0.7600 ;
      RECT 332.5100 0.0000 333.6900 0.7600 ;
      RECT 330.9100 0.0000 332.0900 0.7600 ;
      RECT 329.3100 0.0000 330.4900 0.7600 ;
      RECT 327.7100 0.0000 328.8900 0.7600 ;
      RECT 326.1100 0.0000 327.2900 0.7600 ;
      RECT 324.5100 0.0000 325.6900 0.7600 ;
      RECT 322.9100 0.0000 324.0900 0.7600 ;
      RECT 321.3100 0.0000 322.4900 0.7600 ;
      RECT 319.7100 0.0000 320.8900 0.7600 ;
      RECT 318.1100 0.0000 319.2900 0.7600 ;
      RECT 316.5100 0.0000 317.6900 0.7600 ;
      RECT 314.9100 0.0000 316.0900 0.7600 ;
      RECT 313.3100 0.0000 314.4900 0.7600 ;
      RECT 311.7100 0.0000 312.8900 0.7600 ;
      RECT 310.1100 0.0000 311.2900 0.7600 ;
      RECT 308.5100 0.0000 309.6900 0.7600 ;
      RECT 306.9100 0.0000 308.0900 0.7600 ;
      RECT 305.3100 0.0000 306.4900 0.7600 ;
      RECT 303.7100 0.0000 304.8900 0.7600 ;
      RECT 302.1100 0.0000 303.2900 0.7600 ;
      RECT 300.5100 0.0000 301.6900 0.7600 ;
      RECT 298.9100 0.0000 300.0900 0.7600 ;
      RECT 297.3100 0.0000 298.4900 0.7600 ;
      RECT 295.7100 0.0000 296.8900 0.7600 ;
      RECT 294.1100 0.0000 295.2900 0.7600 ;
      RECT 292.5100 0.0000 293.6900 0.7600 ;
      RECT 290.9100 0.0000 292.0900 0.7600 ;
      RECT 289.3100 0.0000 290.4900 0.7600 ;
      RECT 287.7100 0.0000 288.8900 0.7600 ;
      RECT 286.1100 0.0000 287.2900 0.7600 ;
      RECT 284.5100 0.0000 285.6900 0.7600 ;
      RECT 282.9100 0.0000 284.0900 0.7600 ;
      RECT 281.3100 0.0000 282.4900 0.7600 ;
      RECT 279.7100 0.0000 280.8900 0.7600 ;
      RECT 278.1100 0.0000 279.2900 0.7600 ;
      RECT 276.5100 0.0000 277.6900 0.7600 ;
      RECT 274.9100 0.0000 276.0900 0.7600 ;
      RECT 273.3100 0.0000 274.4900 0.7600 ;
      RECT 271.7100 0.0000 272.8900 0.7600 ;
      RECT 270.1100 0.0000 271.2900 0.7600 ;
      RECT 268.5100 0.0000 269.6900 0.7600 ;
      RECT 266.9100 0.0000 268.0900 0.7600 ;
      RECT 265.3100 0.0000 266.4900 0.7600 ;
      RECT 263.7100 0.0000 264.8900 0.7600 ;
      RECT 262.1100 0.0000 263.2900 0.7600 ;
      RECT 260.5100 0.0000 261.6900 0.7600 ;
      RECT 258.9100 0.0000 260.0900 0.7600 ;
      RECT 257.3100 0.0000 258.4900 0.7600 ;
      RECT 255.7100 0.0000 256.8900 0.7600 ;
      RECT 254.1100 0.0000 255.2900 0.7600 ;
      RECT 252.5100 0.0000 253.6900 0.7600 ;
      RECT 250.9100 0.0000 252.0900 0.7600 ;
      RECT 249.3100 0.0000 250.4900 0.7600 ;
      RECT 247.7100 0.0000 248.8900 0.7600 ;
      RECT 246.1100 0.0000 247.2900 0.7600 ;
      RECT 244.5100 0.0000 245.6900 0.7600 ;
      RECT 242.9100 0.0000 244.0900 0.7600 ;
      RECT 241.3100 0.0000 242.4900 0.7600 ;
      RECT 239.7100 0.0000 240.8900 0.7600 ;
      RECT 238.1100 0.0000 239.2900 0.7600 ;
      RECT 236.5100 0.0000 237.6900 0.7600 ;
      RECT 234.9100 0.0000 236.0900 0.7600 ;
      RECT 233.3100 0.0000 234.4900 0.7600 ;
      RECT 231.7100 0.0000 232.8900 0.7600 ;
      RECT 230.1100 0.0000 231.2900 0.7600 ;
      RECT 228.5100 0.0000 229.6900 0.7600 ;
      RECT 226.9100 0.0000 228.0900 0.7600 ;
      RECT 225.3100 0.0000 226.4900 0.7600 ;
      RECT 223.7100 0.0000 224.8900 0.7600 ;
      RECT 222.1100 0.0000 223.2900 0.7600 ;
      RECT 220.5100 0.0000 221.6900 0.7600 ;
      RECT 218.9100 0.0000 220.0900 0.7600 ;
      RECT 217.3100 0.0000 218.4900 0.7600 ;
      RECT 215.7100 0.0000 216.8900 0.7600 ;
      RECT 214.1100 0.0000 215.2900 0.7600 ;
      RECT 212.5100 0.0000 213.6900 0.7600 ;
      RECT 210.9100 0.0000 212.0900 0.7600 ;
      RECT 209.3100 0.0000 210.4900 0.7600 ;
      RECT 207.7100 0.0000 208.8900 0.7600 ;
      RECT 206.1100 0.0000 207.2900 0.7600 ;
      RECT 204.5100 0.0000 205.6900 0.7600 ;
      RECT 202.9100 0.0000 204.0900 0.7600 ;
      RECT 201.3100 0.0000 202.4900 0.7600 ;
      RECT 199.7100 0.0000 200.8900 0.7600 ;
      RECT 198.1100 0.0000 199.2900 0.7600 ;
      RECT 196.5100 0.0000 197.6900 0.7600 ;
      RECT 194.9100 0.0000 196.0900 0.7600 ;
      RECT 193.3100 0.0000 194.4900 0.7600 ;
      RECT 191.7100 0.0000 192.8900 0.7600 ;
      RECT 190.1100 0.0000 191.2900 0.7600 ;
      RECT 188.5100 0.0000 189.6900 0.7600 ;
      RECT 186.9100 0.0000 188.0900 0.7600 ;
      RECT 185.3100 0.0000 186.4900 0.7600 ;
      RECT 183.7100 0.0000 184.8900 0.7600 ;
      RECT 182.1100 0.0000 183.2900 0.7600 ;
      RECT 180.5100 0.0000 181.6900 0.7600 ;
      RECT 178.9100 0.0000 180.0900 0.7600 ;
      RECT 177.3100 0.0000 178.4900 0.7600 ;
      RECT 175.7100 0.0000 176.8900 0.7600 ;
      RECT 174.1100 0.0000 175.2900 0.7600 ;
      RECT 172.5100 0.0000 173.6900 0.7600 ;
      RECT 170.9100 0.0000 172.0900 0.7600 ;
      RECT 169.3100 0.0000 170.4900 0.7600 ;
      RECT 167.7100 0.0000 168.8900 0.7600 ;
      RECT 166.1100 0.0000 167.2900 0.7600 ;
      RECT 164.5100 0.0000 165.6900 0.7600 ;
      RECT 162.9100 0.0000 164.0900 0.7600 ;
      RECT 161.3100 0.0000 162.4900 0.7600 ;
      RECT 159.7100 0.0000 160.8900 0.7600 ;
      RECT 158.1100 0.0000 159.2900 0.7600 ;
      RECT 156.5100 0.0000 157.6900 0.7600 ;
      RECT 154.9100 0.0000 156.0900 0.7600 ;
      RECT 153.3100 0.0000 154.4900 0.7600 ;
      RECT 151.7100 0.0000 152.8900 0.7600 ;
      RECT 150.1100 0.0000 151.2900 0.7600 ;
      RECT 148.5100 0.0000 149.6900 0.7600 ;
      RECT 146.9100 0.0000 148.0900 0.7600 ;
      RECT 145.3100 0.0000 146.4900 0.7600 ;
      RECT 143.7100 0.0000 144.8900 0.7600 ;
      RECT 142.1100 0.0000 143.2900 0.7600 ;
      RECT 140.5100 0.0000 141.6900 0.7600 ;
      RECT 138.9100 0.0000 140.0900 0.7600 ;
      RECT 137.3100 0.0000 138.4900 0.7600 ;
      RECT 135.7100 0.0000 136.8900 0.7600 ;
      RECT 134.1100 0.0000 135.2900 0.7600 ;
      RECT 132.5100 0.0000 133.6900 0.7600 ;
      RECT 130.9100 0.0000 132.0900 0.7600 ;
      RECT 129.3100 0.0000 130.4900 0.7600 ;
      RECT 127.7100 0.0000 128.8900 0.7600 ;
      RECT 126.1100 0.0000 127.2900 0.7600 ;
      RECT 124.5100 0.0000 125.6900 0.7600 ;
      RECT 122.9100 0.0000 124.0900 0.7600 ;
      RECT 121.3100 0.0000 122.4900 0.7600 ;
      RECT 119.7100 0.0000 120.8900 0.7600 ;
      RECT 118.1100 0.0000 119.2900 0.7600 ;
      RECT 116.5100 0.0000 117.6900 0.7600 ;
      RECT 114.9100 0.0000 116.0900 0.7600 ;
      RECT 113.3100 0.0000 114.4900 0.7600 ;
      RECT 111.7100 0.0000 112.8900 0.7600 ;
      RECT 110.1100 0.0000 111.2900 0.7600 ;
      RECT 108.5100 0.0000 109.6900 0.7600 ;
      RECT 106.9100 0.0000 108.0900 0.7600 ;
      RECT 105.3100 0.0000 106.4900 0.7600 ;
      RECT 103.7100 0.0000 104.8900 0.7600 ;
      RECT 102.1100 0.0000 103.2900 0.7600 ;
      RECT 100.5100 0.0000 101.6900 0.7600 ;
      RECT 98.9100 0.0000 100.0900 0.7600 ;
      RECT 97.3100 0.0000 98.4900 0.7600 ;
      RECT 95.7100 0.0000 96.8900 0.7600 ;
      RECT 94.1100 0.0000 95.2900 0.7600 ;
      RECT 92.5100 0.0000 93.6900 0.7600 ;
      RECT 90.9100 0.0000 92.0900 0.7600 ;
      RECT 89.3100 0.0000 90.4900 0.7600 ;
      RECT 87.7100 0.0000 88.8900 0.7600 ;
      RECT 86.1100 0.0000 87.2900 0.7600 ;
      RECT 84.5100 0.0000 85.6900 0.7600 ;
      RECT 82.9100 0.0000 84.0900 0.7600 ;
      RECT 81.3100 0.0000 82.4900 0.7600 ;
      RECT 79.7100 0.0000 80.8900 0.7600 ;
      RECT 78.1100 0.0000 79.2900 0.7600 ;
      RECT 76.5100 0.0000 77.6900 0.7600 ;
      RECT 74.9100 0.0000 76.0900 0.7600 ;
      RECT 73.3100 0.0000 74.4900 0.7600 ;
      RECT 71.7100 0.0000 72.8900 0.7600 ;
      RECT 70.1100 0.0000 71.2900 0.7600 ;
      RECT 68.5100 0.0000 69.6900 0.7600 ;
      RECT 66.9100 0.0000 68.0900 0.7600 ;
      RECT 65.3100 0.0000 66.4900 0.7600 ;
      RECT 63.7100 0.0000 64.8900 0.7600 ;
      RECT 62.1100 0.0000 63.2900 0.7600 ;
      RECT 60.5100 0.0000 61.6900 0.7600 ;
      RECT 58.9100 0.0000 60.0900 0.7600 ;
      RECT 57.3100 0.0000 58.4900 0.7600 ;
      RECT 55.7100 0.0000 56.8900 0.7600 ;
      RECT 54.1100 0.0000 55.2900 0.7600 ;
      RECT 52.5100 0.0000 53.6900 0.7600 ;
      RECT 50.9100 0.0000 52.0900 0.7600 ;
      RECT 49.3100 0.0000 50.4900 0.7600 ;
      RECT 47.7100 0.0000 48.8900 0.7600 ;
      RECT 46.1100 0.0000 47.2900 0.7600 ;
      RECT 44.5100 0.0000 45.6900 0.7600 ;
      RECT 42.9100 0.0000 44.0900 0.7600 ;
      RECT 41.3100 0.0000 42.4900 0.7600 ;
      RECT 39.7100 0.0000 40.8900 0.7600 ;
      RECT 38.1100 0.0000 39.2900 0.7600 ;
      RECT 36.5100 0.0000 37.6900 0.7600 ;
      RECT 34.9100 0.0000 36.0900 0.7600 ;
      RECT 33.3100 0.0000 34.4900 0.7600 ;
      RECT 31.7100 0.0000 32.8900 0.7600 ;
      RECT 30.1100 0.0000 31.2900 0.7600 ;
      RECT 28.5100 0.0000 29.6900 0.7600 ;
      RECT 26.9100 0.0000 28.0900 0.7600 ;
      RECT 25.3100 0.0000 26.4900 0.7600 ;
      RECT 0.0000 0.0000 24.8900 0.7600 ;
    LAYER M4 ;
      RECT 0.0000 93.4650 450.2000 102.8000 ;
      RECT 293.6300 93.3000 417.6950 93.4650 ;
      RECT 166.5650 93.3000 290.6300 93.4650 ;
      RECT 39.5000 93.3000 163.5650 93.4650 ;
      RECT 0.0000 93.3000 36.5000 93.4650 ;
      RECT 413.6950 9.5000 417.6950 93.3000 ;
      RECT 293.6300 9.5000 410.6950 93.3000 ;
      RECT 286.6300 9.5000 290.6300 93.3000 ;
      RECT 166.5650 9.5000 283.6300 93.3000 ;
      RECT 159.5650 9.5000 163.5650 93.3000 ;
      RECT 39.5000 9.5000 156.5650 93.3000 ;
      RECT 32.5000 9.5000 36.5000 93.3000 ;
      RECT 0.0000 9.5000 29.5000 93.3000 ;
      RECT 420.6950 9.3350 450.2000 93.4650 ;
      RECT 293.6300 9.3350 417.6950 9.5000 ;
      RECT 166.5650 9.3350 290.6300 9.5000 ;
      RECT 39.5000 9.3350 163.5650 9.5000 ;
      RECT 0.0000 9.3350 36.5000 9.5000 ;
      RECT 0.0000 0.0000 450.2000 9.3350 ;
  END
END sram_w16_256

END LIBRARY
