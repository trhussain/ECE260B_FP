##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 22 00:02:49 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 402.4000 BY 401.6000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 0.1500 0.6000 0.2500 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 356.5500 0.6000 356.6500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 352.1500 0.6000 352.2500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 347.7500 0.6000 347.8500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 343.3500 0.6000 343.4500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 338.9500 0.6000 339.0500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 334.5500 0.6000 334.6500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 330.1500 0.6000 330.2500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 325.7500 0.6000 325.8500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 321.3500 0.6000 321.4500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 316.9500 0.6000 317.0500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 312.5500 0.6000 312.6500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 308.1500 0.6000 308.2500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 303.7500 0.6000 303.8500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 299.3500 0.6000 299.4500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 294.9500 0.6000 295.0500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 290.5500 0.6000 290.6500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 286.1500 0.6000 286.2500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 281.7500 0.6000 281.8500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 277.3500 0.6000 277.4500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 272.9500 0.6000 273.0500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 268.5500 0.6000 268.6500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 264.1500 0.6000 264.2500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 259.7500 0.6000 259.8500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 255.3500 0.6000 255.4500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 250.9500 0.6000 251.0500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 246.5500 0.6000 246.6500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 242.1500 0.6000 242.2500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 237.7500 0.6000 237.8500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 233.3500 0.6000 233.4500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 228.9500 0.6000 229.0500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 224.5500 0.6000 224.6500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 220.1500 0.6000 220.2500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 215.7500 0.6000 215.8500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 211.3500 0.6000 211.4500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 206.9500 0.6000 207.0500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 202.5500 0.6000 202.6500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 198.1500 0.6000 198.2500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 193.7500 0.6000 193.8500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 189.3500 0.6000 189.4500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 184.9500 0.6000 185.0500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 180.5500 0.6000 180.6500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 176.1500 0.6000 176.2500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 171.7500 0.6000 171.8500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 167.3500 0.6000 167.4500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 162.9500 0.6000 163.0500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 158.5500 0.6000 158.6500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 154.1500 0.6000 154.2500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 149.7500 0.6000 149.8500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 145.3500 0.6000 145.4500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 140.9500 0.6000 141.0500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 136.5500 0.6000 136.6500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 132.1500 0.6000 132.2500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 127.7500 0.6000 127.8500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 123.3500 0.6000 123.4500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 118.9500 0.6000 119.0500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 114.5500 0.6000 114.6500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 110.1500 0.6000 110.2500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 105.7500 0.6000 105.8500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 101.3500 0.6000 101.4500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 96.9500 0.6000 97.0500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 92.5500 0.6000 92.6500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 88.1500 0.6000 88.2500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 83.7500 0.6000 83.8500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 79.3500 0.6000 79.4500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 19.7500 402.4000 19.8500 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 22.1500 402.4000 22.2500 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 24.5500 402.4000 24.6500 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 26.9500 402.4000 27.0500 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 29.3500 402.4000 29.4500 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 31.7500 402.4000 31.8500 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 34.1500 402.4000 34.2500 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 36.5500 402.4000 36.6500 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 38.9500 402.4000 39.0500 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 41.3500 402.4000 41.4500 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 43.7500 402.4000 43.8500 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 46.1500 402.4000 46.2500 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 48.5500 402.4000 48.6500 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 50.9500 402.4000 51.0500 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 53.3500 402.4000 53.4500 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 55.7500 402.4000 55.8500 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 58.1500 402.4000 58.2500 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 60.5500 402.4000 60.6500 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 62.9500 402.4000 63.0500 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 65.3500 402.4000 65.4500 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 67.7500 402.4000 67.8500 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 70.1500 402.4000 70.2500 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 72.5500 402.4000 72.6500 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 74.9500 402.4000 75.0500 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 77.3500 402.4000 77.4500 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 79.7500 402.4000 79.8500 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 82.1500 402.4000 82.2500 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 84.5500 402.4000 84.6500 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 86.9500 402.4000 87.0500 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 89.3500 402.4000 89.4500 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 91.7500 402.4000 91.8500 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 94.1500 402.4000 94.2500 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 96.5500 402.4000 96.6500 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 98.9500 402.4000 99.0500 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 101.3500 402.4000 101.4500 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 103.7500 402.4000 103.8500 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 106.1500 402.4000 106.2500 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 108.5500 402.4000 108.6500 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 110.9500 402.4000 111.0500 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 113.3500 402.4000 113.4500 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 115.7500 402.4000 115.8500 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 118.1500 402.4000 118.2500 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 120.5500 402.4000 120.6500 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 122.9500 402.4000 123.0500 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 125.3500 402.4000 125.4500 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 127.7500 402.4000 127.8500 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 130.1500 402.4000 130.2500 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 132.5500 402.4000 132.6500 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 134.9500 402.4000 135.0500 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 137.3500 402.4000 137.4500 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 139.7500 402.4000 139.8500 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 142.1500 402.4000 142.2500 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 144.5500 402.4000 144.6500 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 146.9500 402.4000 147.0500 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 149.3500 402.4000 149.4500 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 151.7500 402.4000 151.8500 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 154.1500 402.4000 154.2500 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 156.5500 402.4000 156.6500 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 158.9500 402.4000 159.0500 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 161.3500 402.4000 161.4500 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 163.7500 402.4000 163.8500 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 166.1500 402.4000 166.2500 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 168.5500 402.4000 168.6500 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 170.9500 402.4000 171.0500 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 173.3500 402.4000 173.4500 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 175.7500 402.4000 175.8500 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 178.1500 402.4000 178.2500 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 180.5500 402.4000 180.6500 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 182.9500 402.4000 183.0500 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 185.3500 402.4000 185.4500 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 187.7500 402.4000 187.8500 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 190.1500 402.4000 190.2500 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 192.5500 402.4000 192.6500 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 194.9500 402.4000 195.0500 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 197.3500 402.4000 197.4500 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 199.7500 402.4000 199.8500 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 202.1500 402.4000 202.2500 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 204.5500 402.4000 204.6500 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 206.9500 402.4000 207.0500 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 209.3500 402.4000 209.4500 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 211.7500 402.4000 211.8500 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 214.1500 402.4000 214.2500 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 216.5500 402.4000 216.6500 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 218.9500 402.4000 219.0500 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 221.3500 402.4000 221.4500 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 223.7500 402.4000 223.8500 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 226.1500 402.4000 226.2500 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 228.5500 402.4000 228.6500 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 230.9500 402.4000 231.0500 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 233.3500 402.4000 233.4500 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 235.7500 402.4000 235.8500 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 238.1500 402.4000 238.2500 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 240.5500 402.4000 240.6500 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 242.9500 402.4000 243.0500 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 245.3500 402.4000 245.4500 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 247.7500 402.4000 247.8500 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 250.1500 402.4000 250.2500 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 252.5500 402.4000 252.6500 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 254.9500 402.4000 255.0500 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 257.3500 402.4000 257.4500 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 259.7500 402.4000 259.8500 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 262.1500 402.4000 262.2500 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 264.5500 402.4000 264.6500 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 266.9500 402.4000 267.0500 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 269.3500 402.4000 269.4500 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 271.7500 402.4000 271.8500 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 274.1500 402.4000 274.2500 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 276.5500 402.4000 276.6500 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 278.9500 402.4000 279.0500 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 281.3500 402.4000 281.4500 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 283.7500 402.4000 283.8500 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 286.1500 402.4000 286.2500 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 288.5500 402.4000 288.6500 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 290.9500 402.4000 291.0500 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 293.3500 402.4000 293.4500 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 295.7500 402.4000 295.8500 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 298.1500 402.4000 298.2500 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 300.5500 402.4000 300.6500 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 302.9500 402.4000 303.0500 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 305.3500 402.4000 305.4500 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 307.7500 402.4000 307.8500 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 310.1500 402.4000 310.2500 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 312.5500 402.4000 312.6500 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 314.9500 402.4000 315.0500 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 317.3500 402.4000 317.4500 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 319.7500 402.4000 319.8500 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 322.1500 402.4000 322.2500 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 324.5500 402.4000 324.6500 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 326.9500 402.4000 327.0500 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 329.3500 402.4000 329.4500 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 331.7500 402.4000 331.8500 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 334.1500 402.4000 334.2500 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 336.5500 402.4000 336.6500 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 338.9500 402.4000 339.0500 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 341.3500 402.4000 341.4500 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 343.7500 402.4000 343.8500 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 346.1500 402.4000 346.2500 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 348.5500 402.4000 348.6500 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 350.9500 402.4000 351.0500 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 353.3500 402.4000 353.4500 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 355.7500 402.4000 355.8500 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 358.1500 402.4000 358.2500 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 360.5500 402.4000 360.6500 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 362.9500 402.4000 363.0500 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 365.3500 402.4000 365.4500 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 367.7500 402.4000 367.8500 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 370.1500 402.4000 370.2500 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 372.5500 402.4000 372.6500 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 374.9500 402.4000 375.0500 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 377.3500 402.4000 377.4500 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 379.7500 402.4000 379.8500 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 382.1500 402.4000 382.2500 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 384.5500 402.4000 384.6500 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 386.9500 402.4000 387.0500 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 389.3500 402.4000 389.4500 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 391.7500 402.4000 391.8500 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 394.1500 402.4000 394.2500 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 396.5500 402.4000 396.6500 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 398.9500 402.4000 399.0500 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.8800 401.3500 402.4000 401.4500 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 74.9500 0.6000 75.0500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 70.5500 0.6000 70.6500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 66.1500 0.6000 66.2500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.7500 0.6000 61.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.3500 0.6000 57.4500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 52.9500 0.6000 53.0500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 48.5500 0.6000 48.6500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 44.1500 0.6000 44.2500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 39.7500 0.6000 39.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 35.3500 0.6000 35.4500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.9500 0.6000 31.0500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.5500 0.6000 26.6500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.1500 0.6000 22.2500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.7500 0.6000 17.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 13.3500 0.6000 13.4500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 8.9500 0.6000 9.0500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 4.5500 0.6000 4.6500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 360.9500 0.6000 361.0500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 402.4000 401.6000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 402.4000 401.6000 ;
    LAYER M3 ;
      RECT 0.0000 401.5500 402.4000 401.6000 ;
      RECT 0.0000 401.2500 401.7800 401.5500 ;
      RECT 0.0000 399.1500 402.4000 401.2500 ;
      RECT 0.0000 398.8500 401.7800 399.1500 ;
      RECT 0.0000 396.7500 402.4000 398.8500 ;
      RECT 0.0000 396.4500 401.7800 396.7500 ;
      RECT 0.0000 394.3500 402.4000 396.4500 ;
      RECT 0.0000 394.0500 401.7800 394.3500 ;
      RECT 0.0000 391.9500 402.4000 394.0500 ;
      RECT 0.0000 391.6500 401.7800 391.9500 ;
      RECT 0.0000 389.5500 402.4000 391.6500 ;
      RECT 0.0000 389.2500 401.7800 389.5500 ;
      RECT 0.0000 387.1500 402.4000 389.2500 ;
      RECT 0.0000 386.8500 401.7800 387.1500 ;
      RECT 0.0000 384.7500 402.4000 386.8500 ;
      RECT 0.0000 384.4500 401.7800 384.7500 ;
      RECT 0.0000 382.3500 402.4000 384.4500 ;
      RECT 0.0000 382.0500 401.7800 382.3500 ;
      RECT 0.0000 379.9500 402.4000 382.0500 ;
      RECT 0.0000 379.6500 401.7800 379.9500 ;
      RECT 0.0000 377.5500 402.4000 379.6500 ;
      RECT 0.0000 377.2500 401.7800 377.5500 ;
      RECT 0.0000 375.1500 402.4000 377.2500 ;
      RECT 0.0000 374.8500 401.7800 375.1500 ;
      RECT 0.0000 372.7500 402.4000 374.8500 ;
      RECT 0.0000 372.4500 401.7800 372.7500 ;
      RECT 0.0000 370.3500 402.4000 372.4500 ;
      RECT 0.0000 370.0500 401.7800 370.3500 ;
      RECT 0.0000 367.9500 402.4000 370.0500 ;
      RECT 0.0000 367.6500 401.7800 367.9500 ;
      RECT 0.0000 365.5500 402.4000 367.6500 ;
      RECT 0.0000 365.2500 401.7800 365.5500 ;
      RECT 0.0000 363.1500 402.4000 365.2500 ;
      RECT 0.0000 362.8500 401.7800 363.1500 ;
      RECT 0.0000 361.1500 402.4000 362.8500 ;
      RECT 0.7000 360.8500 402.4000 361.1500 ;
      RECT 0.0000 360.7500 402.4000 360.8500 ;
      RECT 0.0000 360.4500 401.7800 360.7500 ;
      RECT 0.0000 358.3500 402.4000 360.4500 ;
      RECT 0.0000 358.0500 401.7800 358.3500 ;
      RECT 0.0000 356.7500 402.4000 358.0500 ;
      RECT 0.7000 356.4500 402.4000 356.7500 ;
      RECT 0.0000 355.9500 402.4000 356.4500 ;
      RECT 0.0000 355.6500 401.7800 355.9500 ;
      RECT 0.0000 353.5500 402.4000 355.6500 ;
      RECT 0.0000 353.2500 401.7800 353.5500 ;
      RECT 0.0000 352.3500 402.4000 353.2500 ;
      RECT 0.7000 352.0500 402.4000 352.3500 ;
      RECT 0.0000 351.1500 402.4000 352.0500 ;
      RECT 0.0000 350.8500 401.7800 351.1500 ;
      RECT 0.0000 348.7500 402.4000 350.8500 ;
      RECT 0.0000 348.4500 401.7800 348.7500 ;
      RECT 0.0000 347.9500 402.4000 348.4500 ;
      RECT 0.7000 347.6500 402.4000 347.9500 ;
      RECT 0.0000 346.3500 402.4000 347.6500 ;
      RECT 0.0000 346.0500 401.7800 346.3500 ;
      RECT 0.0000 343.9500 402.4000 346.0500 ;
      RECT 0.0000 343.6500 401.7800 343.9500 ;
      RECT 0.0000 343.5500 402.4000 343.6500 ;
      RECT 0.7000 343.2500 402.4000 343.5500 ;
      RECT 0.0000 341.5500 402.4000 343.2500 ;
      RECT 0.0000 341.2500 401.7800 341.5500 ;
      RECT 0.0000 339.1500 402.4000 341.2500 ;
      RECT 0.7000 338.8500 401.7800 339.1500 ;
      RECT 0.0000 336.7500 402.4000 338.8500 ;
      RECT 0.0000 336.4500 401.7800 336.7500 ;
      RECT 0.0000 334.7500 402.4000 336.4500 ;
      RECT 0.7000 334.4500 402.4000 334.7500 ;
      RECT 0.0000 334.3500 402.4000 334.4500 ;
      RECT 0.0000 334.0500 401.7800 334.3500 ;
      RECT 0.0000 331.9500 402.4000 334.0500 ;
      RECT 0.0000 331.6500 401.7800 331.9500 ;
      RECT 0.0000 330.3500 402.4000 331.6500 ;
      RECT 0.7000 330.0500 402.4000 330.3500 ;
      RECT 0.0000 329.5500 402.4000 330.0500 ;
      RECT 0.0000 329.2500 401.7800 329.5500 ;
      RECT 0.0000 327.1500 402.4000 329.2500 ;
      RECT 0.0000 326.8500 401.7800 327.1500 ;
      RECT 0.0000 325.9500 402.4000 326.8500 ;
      RECT 0.7000 325.6500 402.4000 325.9500 ;
      RECT 0.0000 324.7500 402.4000 325.6500 ;
      RECT 0.0000 324.4500 401.7800 324.7500 ;
      RECT 0.0000 322.3500 402.4000 324.4500 ;
      RECT 0.0000 322.0500 401.7800 322.3500 ;
      RECT 0.0000 321.5500 402.4000 322.0500 ;
      RECT 0.7000 321.2500 402.4000 321.5500 ;
      RECT 0.0000 319.9500 402.4000 321.2500 ;
      RECT 0.0000 319.6500 401.7800 319.9500 ;
      RECT 0.0000 317.5500 402.4000 319.6500 ;
      RECT 0.0000 317.2500 401.7800 317.5500 ;
      RECT 0.0000 317.1500 402.4000 317.2500 ;
      RECT 0.7000 316.8500 402.4000 317.1500 ;
      RECT 0.0000 315.1500 402.4000 316.8500 ;
      RECT 0.0000 314.8500 401.7800 315.1500 ;
      RECT 0.0000 312.7500 402.4000 314.8500 ;
      RECT 0.7000 312.4500 401.7800 312.7500 ;
      RECT 0.0000 310.3500 402.4000 312.4500 ;
      RECT 0.0000 310.0500 401.7800 310.3500 ;
      RECT 0.0000 308.3500 402.4000 310.0500 ;
      RECT 0.7000 308.0500 402.4000 308.3500 ;
      RECT 0.0000 307.9500 402.4000 308.0500 ;
      RECT 0.0000 307.6500 401.7800 307.9500 ;
      RECT 0.0000 305.5500 402.4000 307.6500 ;
      RECT 0.0000 305.2500 401.7800 305.5500 ;
      RECT 0.0000 303.9500 402.4000 305.2500 ;
      RECT 0.7000 303.6500 402.4000 303.9500 ;
      RECT 0.0000 303.1500 402.4000 303.6500 ;
      RECT 0.0000 302.8500 401.7800 303.1500 ;
      RECT 0.0000 300.7500 402.4000 302.8500 ;
      RECT 0.0000 300.4500 401.7800 300.7500 ;
      RECT 0.0000 299.5500 402.4000 300.4500 ;
      RECT 0.7000 299.2500 402.4000 299.5500 ;
      RECT 0.0000 298.3500 402.4000 299.2500 ;
      RECT 0.0000 298.0500 401.7800 298.3500 ;
      RECT 0.0000 295.9500 402.4000 298.0500 ;
      RECT 0.0000 295.6500 401.7800 295.9500 ;
      RECT 0.0000 295.1500 402.4000 295.6500 ;
      RECT 0.7000 294.8500 402.4000 295.1500 ;
      RECT 0.0000 293.5500 402.4000 294.8500 ;
      RECT 0.0000 293.2500 401.7800 293.5500 ;
      RECT 0.0000 291.1500 402.4000 293.2500 ;
      RECT 0.0000 290.8500 401.7800 291.1500 ;
      RECT 0.0000 290.7500 402.4000 290.8500 ;
      RECT 0.7000 290.4500 402.4000 290.7500 ;
      RECT 0.0000 288.7500 402.4000 290.4500 ;
      RECT 0.0000 288.4500 401.7800 288.7500 ;
      RECT 0.0000 286.3500 402.4000 288.4500 ;
      RECT 0.7000 286.0500 401.7800 286.3500 ;
      RECT 0.0000 283.9500 402.4000 286.0500 ;
      RECT 0.0000 283.6500 401.7800 283.9500 ;
      RECT 0.0000 281.9500 402.4000 283.6500 ;
      RECT 0.7000 281.6500 402.4000 281.9500 ;
      RECT 0.0000 281.5500 402.4000 281.6500 ;
      RECT 0.0000 281.2500 401.7800 281.5500 ;
      RECT 0.0000 279.1500 402.4000 281.2500 ;
      RECT 0.0000 278.8500 401.7800 279.1500 ;
      RECT 0.0000 277.5500 402.4000 278.8500 ;
      RECT 0.7000 277.2500 402.4000 277.5500 ;
      RECT 0.0000 276.7500 402.4000 277.2500 ;
      RECT 0.0000 276.4500 401.7800 276.7500 ;
      RECT 0.0000 274.3500 402.4000 276.4500 ;
      RECT 0.0000 274.0500 401.7800 274.3500 ;
      RECT 0.0000 273.1500 402.4000 274.0500 ;
      RECT 0.7000 272.8500 402.4000 273.1500 ;
      RECT 0.0000 271.9500 402.4000 272.8500 ;
      RECT 0.0000 271.6500 401.7800 271.9500 ;
      RECT 0.0000 269.5500 402.4000 271.6500 ;
      RECT 0.0000 269.2500 401.7800 269.5500 ;
      RECT 0.0000 268.7500 402.4000 269.2500 ;
      RECT 0.7000 268.4500 402.4000 268.7500 ;
      RECT 0.0000 267.1500 402.4000 268.4500 ;
      RECT 0.0000 266.8500 401.7800 267.1500 ;
      RECT 0.0000 264.7500 402.4000 266.8500 ;
      RECT 0.0000 264.4500 401.7800 264.7500 ;
      RECT 0.0000 264.3500 402.4000 264.4500 ;
      RECT 0.7000 264.0500 402.4000 264.3500 ;
      RECT 0.0000 262.3500 402.4000 264.0500 ;
      RECT 0.0000 262.0500 401.7800 262.3500 ;
      RECT 0.0000 259.9500 402.4000 262.0500 ;
      RECT 0.7000 259.6500 401.7800 259.9500 ;
      RECT 0.0000 257.5500 402.4000 259.6500 ;
      RECT 0.0000 257.2500 401.7800 257.5500 ;
      RECT 0.0000 255.5500 402.4000 257.2500 ;
      RECT 0.7000 255.2500 402.4000 255.5500 ;
      RECT 0.0000 255.1500 402.4000 255.2500 ;
      RECT 0.0000 254.8500 401.7800 255.1500 ;
      RECT 0.0000 252.7500 402.4000 254.8500 ;
      RECT 0.0000 252.4500 401.7800 252.7500 ;
      RECT 0.0000 251.1500 402.4000 252.4500 ;
      RECT 0.7000 250.8500 402.4000 251.1500 ;
      RECT 0.0000 250.3500 402.4000 250.8500 ;
      RECT 0.0000 250.0500 401.7800 250.3500 ;
      RECT 0.0000 247.9500 402.4000 250.0500 ;
      RECT 0.0000 247.6500 401.7800 247.9500 ;
      RECT 0.0000 246.7500 402.4000 247.6500 ;
      RECT 0.7000 246.4500 402.4000 246.7500 ;
      RECT 0.0000 245.5500 402.4000 246.4500 ;
      RECT 0.0000 245.2500 401.7800 245.5500 ;
      RECT 0.0000 243.1500 402.4000 245.2500 ;
      RECT 0.0000 242.8500 401.7800 243.1500 ;
      RECT 0.0000 242.3500 402.4000 242.8500 ;
      RECT 0.7000 242.0500 402.4000 242.3500 ;
      RECT 0.0000 240.7500 402.4000 242.0500 ;
      RECT 0.0000 240.4500 401.7800 240.7500 ;
      RECT 0.0000 238.3500 402.4000 240.4500 ;
      RECT 0.0000 238.0500 401.7800 238.3500 ;
      RECT 0.0000 237.9500 402.4000 238.0500 ;
      RECT 0.7000 237.6500 402.4000 237.9500 ;
      RECT 0.0000 235.9500 402.4000 237.6500 ;
      RECT 0.0000 235.6500 401.7800 235.9500 ;
      RECT 0.0000 233.5500 402.4000 235.6500 ;
      RECT 0.7000 233.2500 401.7800 233.5500 ;
      RECT 0.0000 231.1500 402.4000 233.2500 ;
      RECT 0.0000 230.8500 401.7800 231.1500 ;
      RECT 0.0000 229.1500 402.4000 230.8500 ;
      RECT 0.7000 228.8500 402.4000 229.1500 ;
      RECT 0.0000 228.7500 402.4000 228.8500 ;
      RECT 0.0000 228.4500 401.7800 228.7500 ;
      RECT 0.0000 226.3500 402.4000 228.4500 ;
      RECT 0.0000 226.0500 401.7800 226.3500 ;
      RECT 0.0000 224.7500 402.4000 226.0500 ;
      RECT 0.7000 224.4500 402.4000 224.7500 ;
      RECT 0.0000 223.9500 402.4000 224.4500 ;
      RECT 0.0000 223.6500 401.7800 223.9500 ;
      RECT 0.0000 221.5500 402.4000 223.6500 ;
      RECT 0.0000 221.2500 401.7800 221.5500 ;
      RECT 0.0000 220.3500 402.4000 221.2500 ;
      RECT 0.7000 220.0500 402.4000 220.3500 ;
      RECT 0.0000 219.1500 402.4000 220.0500 ;
      RECT 0.0000 218.8500 401.7800 219.1500 ;
      RECT 0.0000 216.7500 402.4000 218.8500 ;
      RECT 0.0000 216.4500 401.7800 216.7500 ;
      RECT 0.0000 215.9500 402.4000 216.4500 ;
      RECT 0.7000 215.6500 402.4000 215.9500 ;
      RECT 0.0000 214.3500 402.4000 215.6500 ;
      RECT 0.0000 214.0500 401.7800 214.3500 ;
      RECT 0.0000 211.9500 402.4000 214.0500 ;
      RECT 0.0000 211.6500 401.7800 211.9500 ;
      RECT 0.0000 211.5500 402.4000 211.6500 ;
      RECT 0.7000 211.2500 402.4000 211.5500 ;
      RECT 0.0000 209.5500 402.4000 211.2500 ;
      RECT 0.0000 209.2500 401.7800 209.5500 ;
      RECT 0.0000 207.1500 402.4000 209.2500 ;
      RECT 0.7000 206.8500 401.7800 207.1500 ;
      RECT 0.0000 204.7500 402.4000 206.8500 ;
      RECT 0.0000 204.4500 401.7800 204.7500 ;
      RECT 0.0000 202.7500 402.4000 204.4500 ;
      RECT 0.7000 202.4500 402.4000 202.7500 ;
      RECT 0.0000 202.3500 402.4000 202.4500 ;
      RECT 0.0000 202.0500 401.7800 202.3500 ;
      RECT 0.0000 199.9500 402.4000 202.0500 ;
      RECT 0.0000 199.6500 401.7800 199.9500 ;
      RECT 0.0000 198.3500 402.4000 199.6500 ;
      RECT 0.7000 198.0500 402.4000 198.3500 ;
      RECT 0.0000 197.5500 402.4000 198.0500 ;
      RECT 0.0000 197.2500 401.7800 197.5500 ;
      RECT 0.0000 195.1500 402.4000 197.2500 ;
      RECT 0.0000 194.8500 401.7800 195.1500 ;
      RECT 0.0000 193.9500 402.4000 194.8500 ;
      RECT 0.7000 193.6500 402.4000 193.9500 ;
      RECT 0.0000 192.7500 402.4000 193.6500 ;
      RECT 0.0000 192.4500 401.7800 192.7500 ;
      RECT 0.0000 190.3500 402.4000 192.4500 ;
      RECT 0.0000 190.0500 401.7800 190.3500 ;
      RECT 0.0000 189.5500 402.4000 190.0500 ;
      RECT 0.7000 189.2500 402.4000 189.5500 ;
      RECT 0.0000 187.9500 402.4000 189.2500 ;
      RECT 0.0000 187.6500 401.7800 187.9500 ;
      RECT 0.0000 185.5500 402.4000 187.6500 ;
      RECT 0.0000 185.2500 401.7800 185.5500 ;
      RECT 0.0000 185.1500 402.4000 185.2500 ;
      RECT 0.7000 184.8500 402.4000 185.1500 ;
      RECT 0.0000 183.1500 402.4000 184.8500 ;
      RECT 0.0000 182.8500 401.7800 183.1500 ;
      RECT 0.0000 180.7500 402.4000 182.8500 ;
      RECT 0.7000 180.4500 401.7800 180.7500 ;
      RECT 0.0000 178.3500 402.4000 180.4500 ;
      RECT 0.0000 178.0500 401.7800 178.3500 ;
      RECT 0.0000 176.3500 402.4000 178.0500 ;
      RECT 0.7000 176.0500 402.4000 176.3500 ;
      RECT 0.0000 175.9500 402.4000 176.0500 ;
      RECT 0.0000 175.6500 401.7800 175.9500 ;
      RECT 0.0000 173.5500 402.4000 175.6500 ;
      RECT 0.0000 173.2500 401.7800 173.5500 ;
      RECT 0.0000 171.9500 402.4000 173.2500 ;
      RECT 0.7000 171.6500 402.4000 171.9500 ;
      RECT 0.0000 171.1500 402.4000 171.6500 ;
      RECT 0.0000 170.8500 401.7800 171.1500 ;
      RECT 0.0000 168.7500 402.4000 170.8500 ;
      RECT 0.0000 168.4500 401.7800 168.7500 ;
      RECT 0.0000 167.5500 402.4000 168.4500 ;
      RECT 0.7000 167.2500 402.4000 167.5500 ;
      RECT 0.0000 166.3500 402.4000 167.2500 ;
      RECT 0.0000 166.0500 401.7800 166.3500 ;
      RECT 0.0000 163.9500 402.4000 166.0500 ;
      RECT 0.0000 163.6500 401.7800 163.9500 ;
      RECT 0.0000 163.1500 402.4000 163.6500 ;
      RECT 0.7000 162.8500 402.4000 163.1500 ;
      RECT 0.0000 161.5500 402.4000 162.8500 ;
      RECT 0.0000 161.2500 401.7800 161.5500 ;
      RECT 0.0000 159.1500 402.4000 161.2500 ;
      RECT 0.0000 158.8500 401.7800 159.1500 ;
      RECT 0.0000 158.7500 402.4000 158.8500 ;
      RECT 0.7000 158.4500 402.4000 158.7500 ;
      RECT 0.0000 156.7500 402.4000 158.4500 ;
      RECT 0.0000 156.4500 401.7800 156.7500 ;
      RECT 0.0000 154.3500 402.4000 156.4500 ;
      RECT 0.7000 154.0500 401.7800 154.3500 ;
      RECT 0.0000 151.9500 402.4000 154.0500 ;
      RECT 0.0000 151.6500 401.7800 151.9500 ;
      RECT 0.0000 149.9500 402.4000 151.6500 ;
      RECT 0.7000 149.6500 402.4000 149.9500 ;
      RECT 0.0000 149.5500 402.4000 149.6500 ;
      RECT 0.0000 149.2500 401.7800 149.5500 ;
      RECT 0.0000 147.1500 402.4000 149.2500 ;
      RECT 0.0000 146.8500 401.7800 147.1500 ;
      RECT 0.0000 145.5500 402.4000 146.8500 ;
      RECT 0.7000 145.2500 402.4000 145.5500 ;
      RECT 0.0000 144.7500 402.4000 145.2500 ;
      RECT 0.0000 144.4500 401.7800 144.7500 ;
      RECT 0.0000 142.3500 402.4000 144.4500 ;
      RECT 0.0000 142.0500 401.7800 142.3500 ;
      RECT 0.0000 141.1500 402.4000 142.0500 ;
      RECT 0.7000 140.8500 402.4000 141.1500 ;
      RECT 0.0000 139.9500 402.4000 140.8500 ;
      RECT 0.0000 139.6500 401.7800 139.9500 ;
      RECT 0.0000 137.5500 402.4000 139.6500 ;
      RECT 0.0000 137.2500 401.7800 137.5500 ;
      RECT 0.0000 136.7500 402.4000 137.2500 ;
      RECT 0.7000 136.4500 402.4000 136.7500 ;
      RECT 0.0000 135.1500 402.4000 136.4500 ;
      RECT 0.0000 134.8500 401.7800 135.1500 ;
      RECT 0.0000 132.7500 402.4000 134.8500 ;
      RECT 0.0000 132.4500 401.7800 132.7500 ;
      RECT 0.0000 132.3500 402.4000 132.4500 ;
      RECT 0.7000 132.0500 402.4000 132.3500 ;
      RECT 0.0000 130.3500 402.4000 132.0500 ;
      RECT 0.0000 130.0500 401.7800 130.3500 ;
      RECT 0.0000 127.9500 402.4000 130.0500 ;
      RECT 0.7000 127.6500 401.7800 127.9500 ;
      RECT 0.0000 125.5500 402.4000 127.6500 ;
      RECT 0.0000 125.2500 401.7800 125.5500 ;
      RECT 0.0000 123.5500 402.4000 125.2500 ;
      RECT 0.7000 123.2500 402.4000 123.5500 ;
      RECT 0.0000 123.1500 402.4000 123.2500 ;
      RECT 0.0000 122.8500 401.7800 123.1500 ;
      RECT 0.0000 120.7500 402.4000 122.8500 ;
      RECT 0.0000 120.4500 401.7800 120.7500 ;
      RECT 0.0000 119.1500 402.4000 120.4500 ;
      RECT 0.7000 118.8500 402.4000 119.1500 ;
      RECT 0.0000 118.3500 402.4000 118.8500 ;
      RECT 0.0000 118.0500 401.7800 118.3500 ;
      RECT 0.0000 115.9500 402.4000 118.0500 ;
      RECT 0.0000 115.6500 401.7800 115.9500 ;
      RECT 0.0000 114.7500 402.4000 115.6500 ;
      RECT 0.7000 114.4500 402.4000 114.7500 ;
      RECT 0.0000 113.5500 402.4000 114.4500 ;
      RECT 0.0000 113.2500 401.7800 113.5500 ;
      RECT 0.0000 111.1500 402.4000 113.2500 ;
      RECT 0.0000 110.8500 401.7800 111.1500 ;
      RECT 0.0000 110.3500 402.4000 110.8500 ;
      RECT 0.7000 110.0500 402.4000 110.3500 ;
      RECT 0.0000 108.7500 402.4000 110.0500 ;
      RECT 0.0000 108.4500 401.7800 108.7500 ;
      RECT 0.0000 106.3500 402.4000 108.4500 ;
      RECT 0.0000 106.0500 401.7800 106.3500 ;
      RECT 0.0000 105.9500 402.4000 106.0500 ;
      RECT 0.7000 105.6500 402.4000 105.9500 ;
      RECT 0.0000 103.9500 402.4000 105.6500 ;
      RECT 0.0000 103.6500 401.7800 103.9500 ;
      RECT 0.0000 101.5500 402.4000 103.6500 ;
      RECT 0.7000 101.2500 401.7800 101.5500 ;
      RECT 0.0000 99.1500 402.4000 101.2500 ;
      RECT 0.0000 98.8500 401.7800 99.1500 ;
      RECT 0.0000 97.1500 402.4000 98.8500 ;
      RECT 0.7000 96.8500 402.4000 97.1500 ;
      RECT 0.0000 96.7500 402.4000 96.8500 ;
      RECT 0.0000 96.4500 401.7800 96.7500 ;
      RECT 0.0000 94.3500 402.4000 96.4500 ;
      RECT 0.0000 94.0500 401.7800 94.3500 ;
      RECT 0.0000 92.7500 402.4000 94.0500 ;
      RECT 0.7000 92.4500 402.4000 92.7500 ;
      RECT 0.0000 91.9500 402.4000 92.4500 ;
      RECT 0.0000 91.6500 401.7800 91.9500 ;
      RECT 0.0000 89.5500 402.4000 91.6500 ;
      RECT 0.0000 89.2500 401.7800 89.5500 ;
      RECT 0.0000 88.3500 402.4000 89.2500 ;
      RECT 0.7000 88.0500 402.4000 88.3500 ;
      RECT 0.0000 87.1500 402.4000 88.0500 ;
      RECT 0.0000 86.8500 401.7800 87.1500 ;
      RECT 0.0000 84.7500 402.4000 86.8500 ;
      RECT 0.0000 84.4500 401.7800 84.7500 ;
      RECT 0.0000 83.9500 402.4000 84.4500 ;
      RECT 0.7000 83.6500 402.4000 83.9500 ;
      RECT 0.0000 82.3500 402.4000 83.6500 ;
      RECT 0.0000 82.0500 401.7800 82.3500 ;
      RECT 0.0000 79.9500 402.4000 82.0500 ;
      RECT 0.0000 79.6500 401.7800 79.9500 ;
      RECT 0.0000 79.5500 402.4000 79.6500 ;
      RECT 0.7000 79.2500 402.4000 79.5500 ;
      RECT 0.0000 77.5500 402.4000 79.2500 ;
      RECT 0.0000 77.2500 401.7800 77.5500 ;
      RECT 0.0000 75.1500 402.4000 77.2500 ;
      RECT 0.7000 74.8500 401.7800 75.1500 ;
      RECT 0.0000 72.7500 402.4000 74.8500 ;
      RECT 0.0000 72.4500 401.7800 72.7500 ;
      RECT 0.0000 70.7500 402.4000 72.4500 ;
      RECT 0.7000 70.4500 402.4000 70.7500 ;
      RECT 0.0000 70.3500 402.4000 70.4500 ;
      RECT 0.0000 70.0500 401.7800 70.3500 ;
      RECT 0.0000 67.9500 402.4000 70.0500 ;
      RECT 0.0000 67.6500 401.7800 67.9500 ;
      RECT 0.0000 66.3500 402.4000 67.6500 ;
      RECT 0.7000 66.0500 402.4000 66.3500 ;
      RECT 0.0000 65.5500 402.4000 66.0500 ;
      RECT 0.0000 65.2500 401.7800 65.5500 ;
      RECT 0.0000 63.1500 402.4000 65.2500 ;
      RECT 0.0000 62.8500 401.7800 63.1500 ;
      RECT 0.0000 61.9500 402.4000 62.8500 ;
      RECT 0.7000 61.6500 402.4000 61.9500 ;
      RECT 0.0000 60.7500 402.4000 61.6500 ;
      RECT 0.0000 60.4500 401.7800 60.7500 ;
      RECT 0.0000 58.3500 402.4000 60.4500 ;
      RECT 0.0000 58.0500 401.7800 58.3500 ;
      RECT 0.0000 57.5500 402.4000 58.0500 ;
      RECT 0.7000 57.2500 402.4000 57.5500 ;
      RECT 0.0000 55.9500 402.4000 57.2500 ;
      RECT 0.0000 55.6500 401.7800 55.9500 ;
      RECT 0.0000 53.5500 402.4000 55.6500 ;
      RECT 0.0000 53.2500 401.7800 53.5500 ;
      RECT 0.0000 53.1500 402.4000 53.2500 ;
      RECT 0.7000 52.8500 402.4000 53.1500 ;
      RECT 0.0000 51.1500 402.4000 52.8500 ;
      RECT 0.0000 50.8500 401.7800 51.1500 ;
      RECT 0.0000 48.7500 402.4000 50.8500 ;
      RECT 0.7000 48.4500 401.7800 48.7500 ;
      RECT 0.0000 46.3500 402.4000 48.4500 ;
      RECT 0.0000 46.0500 401.7800 46.3500 ;
      RECT 0.0000 44.3500 402.4000 46.0500 ;
      RECT 0.7000 44.0500 402.4000 44.3500 ;
      RECT 0.0000 43.9500 402.4000 44.0500 ;
      RECT 0.0000 43.6500 401.7800 43.9500 ;
      RECT 0.0000 41.5500 402.4000 43.6500 ;
      RECT 0.0000 41.2500 401.7800 41.5500 ;
      RECT 0.0000 39.9500 402.4000 41.2500 ;
      RECT 0.7000 39.6500 402.4000 39.9500 ;
      RECT 0.0000 39.1500 402.4000 39.6500 ;
      RECT 0.0000 38.8500 401.7800 39.1500 ;
      RECT 0.0000 36.7500 402.4000 38.8500 ;
      RECT 0.0000 36.4500 401.7800 36.7500 ;
      RECT 0.0000 35.5500 402.4000 36.4500 ;
      RECT 0.7000 35.2500 402.4000 35.5500 ;
      RECT 0.0000 34.3500 402.4000 35.2500 ;
      RECT 0.0000 34.0500 401.7800 34.3500 ;
      RECT 0.0000 31.9500 402.4000 34.0500 ;
      RECT 0.0000 31.6500 401.7800 31.9500 ;
      RECT 0.0000 31.1500 402.4000 31.6500 ;
      RECT 0.7000 30.8500 402.4000 31.1500 ;
      RECT 0.0000 29.5500 402.4000 30.8500 ;
      RECT 0.0000 29.2500 401.7800 29.5500 ;
      RECT 0.0000 27.1500 402.4000 29.2500 ;
      RECT 0.0000 26.8500 401.7800 27.1500 ;
      RECT 0.0000 26.7500 402.4000 26.8500 ;
      RECT 0.7000 26.4500 402.4000 26.7500 ;
      RECT 0.0000 24.7500 402.4000 26.4500 ;
      RECT 0.0000 24.4500 401.7800 24.7500 ;
      RECT 0.0000 22.3500 402.4000 24.4500 ;
      RECT 0.7000 22.0500 401.7800 22.3500 ;
      RECT 0.0000 19.9500 402.4000 22.0500 ;
      RECT 0.0000 19.6500 401.7800 19.9500 ;
      RECT 0.0000 17.9500 402.4000 19.6500 ;
      RECT 0.7000 17.6500 402.4000 17.9500 ;
      RECT 0.0000 13.5500 402.4000 17.6500 ;
      RECT 0.7000 13.2500 402.4000 13.5500 ;
      RECT 0.0000 9.1500 402.4000 13.2500 ;
      RECT 0.7000 8.8500 402.4000 9.1500 ;
      RECT 0.0000 4.7500 402.4000 8.8500 ;
      RECT 0.7000 4.4500 402.4000 4.7500 ;
      RECT 0.0000 0.3500 402.4000 4.4500 ;
      RECT 0.7000 0.0500 402.4000 0.3500 ;
      RECT 0.0000 0.0000 402.4000 0.0500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 402.4000 401.6000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 402.4000 401.6000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 402.4000 401.6000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 402.4000 401.6000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 402.4000 401.6000 ;
  END
END core

END LIBRARY
