##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 09:05:40 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16
  CLASS BLOCK ;
  SIZE 268.0000 BY 92.0000 ;
  FOREIGN sram_w16 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 38.1500 0.6000 38.2500 ;
    END
  END CLK
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 228.2500 0.0000 228.3500 0.6000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 226.6500 0.0000 226.7500 0.6000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 225.0500 0.0000 225.1500 0.6000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 223.4500 0.0000 223.5500 0.6000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 221.8500 0.0000 221.9500 0.6000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220.2500 0.0000 220.3500 0.6000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 218.6500 0.0000 218.7500 0.6000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 217.0500 0.0000 217.1500 0.6000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 215.4500 0.0000 215.5500 0.6000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 213.8500 0.0000 213.9500 0.6000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 212.2500 0.0000 212.3500 0.6000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 210.6500 0.0000 210.7500 0.6000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 209.0500 0.0000 209.1500 0.6000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 207.4500 0.0000 207.5500 0.6000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 205.8500 0.0000 205.9500 0.6000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 204.2500 0.0000 204.3500 0.6000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 202.6500 0.0000 202.7500 0.6000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 201.0500 0.0000 201.1500 0.6000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 199.4500 0.0000 199.5500 0.6000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 197.8500 0.0000 197.9500 0.6000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 196.2500 0.0000 196.3500 0.6000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 194.6500 0.0000 194.7500 0.6000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 193.0500 0.0000 193.1500 0.6000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 191.4500 0.0000 191.5500 0.6000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 189.8500 0.0000 189.9500 0.6000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 188.2500 0.0000 188.3500 0.6000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 186.6500 0.0000 186.7500 0.6000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 185.0500 0.0000 185.1500 0.6000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.4500 0.0000 183.5500 0.6000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 181.8500 0.0000 181.9500 0.6000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.2500 0.0000 180.3500 0.6000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.6500 0.0000 178.7500 0.6000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.0500 0.0000 177.1500 0.6000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.4500 0.0000 175.5500 0.6000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.8500 0.0000 173.9500 0.6000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.2500 0.0000 172.3500 0.6000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 170.6500 0.0000 170.7500 0.6000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 169.0500 0.0000 169.1500 0.6000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.4500 0.0000 167.5500 0.6000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.8500 0.0000 165.9500 0.6000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.2500 0.0000 164.3500 0.6000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.6500 0.0000 162.7500 0.6000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.0500 0.0000 161.1500 0.6000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.4500 0.0000 159.5500 0.6000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 157.8500 0.0000 157.9500 0.6000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.2500 0.0000 156.3500 0.6000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.6500 0.0000 154.7500 0.6000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.0500 0.0000 153.1500 0.6000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.4500 0.0000 151.5500 0.6000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 149.8500 0.0000 149.9500 0.6000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.2500 0.0000 148.3500 0.6000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 146.6500 0.0000 146.7500 0.6000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 145.0500 0.0000 145.1500 0.6000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.4500 0.0000 143.5500 0.6000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.8500 0.0000 141.9500 0.6000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.2500 0.0000 140.3500 0.6000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.6500 0.0000 138.7500 0.6000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 137.0500 0.0000 137.1500 0.6000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.4500 0.0000 135.5500 0.6000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 133.8500 0.0000 133.9500 0.6000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.2500 0.0000 132.3500 0.6000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 130.6500 0.0000 130.7500 0.6000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.0500 0.0000 129.1500 0.6000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 127.4500 0.0000 127.5500 0.6000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.8500 0.0000 125.9500 0.6000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.2500 0.0000 124.3500 0.6000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.6500 0.0000 122.7500 0.6000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.0500 0.0000 121.1500 0.6000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.4500 0.0000 119.5500 0.6000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.8500 0.0000 117.9500 0.6000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.2500 0.0000 116.3500 0.6000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.6500 0.0000 114.7500 0.6000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.0500 0.0000 113.1500 0.6000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.4500 0.0000 111.5500 0.6000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.8500 0.0000 109.9500 0.6000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.2500 0.0000 108.3500 0.6000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.6500 0.0000 106.7500 0.6000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.0500 0.0000 105.1500 0.6000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.4500 0.0000 103.5500 0.6000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.8500 0.0000 101.9500 0.6000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.2500 0.0000 100.3500 0.6000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.6500 0.0000 98.7500 0.6000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.0500 0.0000 97.1500 0.6000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.4500 0.0000 95.5500 0.6000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.8500 0.0000 93.9500 0.6000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.2500 0.0000 92.3500 0.6000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.6500 0.0000 90.7500 0.6000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.0500 0.0000 89.1500 0.6000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.4500 0.0000 87.5500 0.6000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.8500 0.0000 85.9500 0.6000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.2500 0.0000 84.3500 0.6000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.6500 0.0000 82.7500 0.6000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.0500 0.0000 81.1500 0.6000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.4500 0.0000 79.5500 0.6000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 77.8500 0.0000 77.9500 0.6000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.2500 0.0000 76.3500 0.6000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 74.6500 0.0000 74.7500 0.6000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.0500 0.0000 73.1500 0.6000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.4500 0.0000 71.5500 0.6000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 69.8500 0.0000 69.9500 0.6000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.2500 0.0000 68.3500 0.6000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 66.6500 0.0000 66.7500 0.6000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.0500 0.0000 65.1500 0.6000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 63.4500 0.0000 63.5500 0.6000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 61.8500 0.0000 61.9500 0.6000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60.2500 0.0000 60.3500 0.6000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.6500 0.0000 58.7500 0.6000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 57.0500 0.0000 57.1500 0.6000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.4500 0.0000 55.5500 0.6000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 53.8500 0.0000 53.9500 0.6000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.2500 0.0000 52.3500 0.6000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 50.6500 0.0000 50.7500 0.6000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 49.0500 0.0000 49.1500 0.6000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 47.4500 0.0000 47.5500 0.6000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 45.8500 0.0000 45.9500 0.6000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 44.2500 0.0000 44.3500 0.6000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 42.6500 0.0000 42.7500 0.6000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 41.0500 0.0000 41.1500 0.6000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.4500 0.0000 39.5500 0.6000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 37.8500 0.0000 37.9500 0.6000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 36.2500 0.0000 36.3500 0.6000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 34.6500 0.0000 34.7500 0.6000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 33.0500 0.0000 33.1500 0.6000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 31.4500 0.0000 31.5500 0.6000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 29.8500 0.0000 29.9500 0.6000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 28.2500 0.0000 28.3500 0.6000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 26.6500 0.0000 26.7500 0.6000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 25.0500 0.0000 25.1500 0.6000 ;
    END
  END D[0]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 228.2500 91.4000 228.3500 92.0000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 226.6500 91.4000 226.7500 92.0000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 225.0500 91.4000 225.1500 92.0000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 223.4500 91.4000 223.5500 92.0000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 221.8500 91.4000 221.9500 92.0000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220.2500 91.4000 220.3500 92.0000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 218.6500 91.4000 218.7500 92.0000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 217.0500 91.4000 217.1500 92.0000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 215.4500 91.4000 215.5500 92.0000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 213.8500 91.4000 213.9500 92.0000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 212.2500 91.4000 212.3500 92.0000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 210.6500 91.4000 210.7500 92.0000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 209.0500 91.4000 209.1500 92.0000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 207.4500 91.4000 207.5500 92.0000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 205.8500 91.4000 205.9500 92.0000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 204.2500 91.4000 204.3500 92.0000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 202.6500 91.4000 202.7500 92.0000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 201.0500 91.4000 201.1500 92.0000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 199.4500 91.4000 199.5500 92.0000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 197.8500 91.4000 197.9500 92.0000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 196.2500 91.4000 196.3500 92.0000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 194.6500 91.4000 194.7500 92.0000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 193.0500 91.4000 193.1500 92.0000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 191.4500 91.4000 191.5500 92.0000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 189.8500 91.4000 189.9500 92.0000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 188.2500 91.4000 188.3500 92.0000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 186.6500 91.4000 186.7500 92.0000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 185.0500 91.4000 185.1500 92.0000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.4500 91.4000 183.5500 92.0000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 181.8500 91.4000 181.9500 92.0000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.2500 91.4000 180.3500 92.0000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.6500 91.4000 178.7500 92.0000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.0500 91.4000 177.1500 92.0000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.4500 91.4000 175.5500 92.0000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.8500 91.4000 173.9500 92.0000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.2500 91.4000 172.3500 92.0000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 170.6500 91.4000 170.7500 92.0000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 169.0500 91.4000 169.1500 92.0000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.4500 91.4000 167.5500 92.0000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.8500 91.4000 165.9500 92.0000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.2500 91.4000 164.3500 92.0000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.6500 91.4000 162.7500 92.0000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.0500 91.4000 161.1500 92.0000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.4500 91.4000 159.5500 92.0000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 157.8500 91.4000 157.9500 92.0000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.2500 91.4000 156.3500 92.0000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.6500 91.4000 154.7500 92.0000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.0500 91.4000 153.1500 92.0000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.4500 91.4000 151.5500 92.0000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 149.8500 91.4000 149.9500 92.0000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.2500 91.4000 148.3500 92.0000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 146.6500 91.4000 146.7500 92.0000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 145.0500 91.4000 145.1500 92.0000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.4500 91.4000 143.5500 92.0000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.8500 91.4000 141.9500 92.0000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.2500 91.4000 140.3500 92.0000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.6500 91.4000 138.7500 92.0000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 137.0500 91.4000 137.1500 92.0000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.4500 91.4000 135.5500 92.0000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 133.8500 91.4000 133.9500 92.0000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.2500 91.4000 132.3500 92.0000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 130.6500 91.4000 130.7500 92.0000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.0500 91.4000 129.1500 92.0000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 127.4500 91.4000 127.5500 92.0000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.8500 91.4000 125.9500 92.0000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.2500 91.4000 124.3500 92.0000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.6500 91.4000 122.7500 92.0000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.0500 91.4000 121.1500 92.0000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.4500 91.4000 119.5500 92.0000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.8500 91.4000 117.9500 92.0000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.2500 91.4000 116.3500 92.0000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.6500 91.4000 114.7500 92.0000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.0500 91.4000 113.1500 92.0000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.4500 91.4000 111.5500 92.0000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.8500 91.4000 109.9500 92.0000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.2500 91.4000 108.3500 92.0000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.6500 91.4000 106.7500 92.0000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.0500 91.4000 105.1500 92.0000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.4500 91.4000 103.5500 92.0000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.8500 91.4000 101.9500 92.0000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.2500 91.4000 100.3500 92.0000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.6500 91.4000 98.7500 92.0000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.0500 91.4000 97.1500 92.0000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.4500 91.4000 95.5500 92.0000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.8500 91.4000 93.9500 92.0000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.2500 91.4000 92.3500 92.0000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.6500 91.4000 90.7500 92.0000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.0500 91.4000 89.1500 92.0000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.4500 91.4000 87.5500 92.0000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.8500 91.4000 85.9500 92.0000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.2500 91.4000 84.3500 92.0000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.6500 91.4000 82.7500 92.0000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.0500 91.4000 81.1500 92.0000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.4500 91.4000 79.5500 92.0000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 77.8500 91.4000 77.9500 92.0000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.2500 91.4000 76.3500 92.0000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 74.6500 91.4000 74.7500 92.0000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.0500 91.4000 73.1500 92.0000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.4500 91.4000 71.5500 92.0000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 69.8500 91.4000 69.9500 92.0000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.2500 91.4000 68.3500 92.0000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 66.6500 91.4000 66.7500 92.0000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.0500 91.4000 65.1500 92.0000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 63.4500 91.4000 63.5500 92.0000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 61.8500 91.4000 61.9500 92.0000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60.2500 91.4000 60.3500 92.0000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.6500 91.4000 58.7500 92.0000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 57.0500 91.4000 57.1500 92.0000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.4500 91.4000 55.5500 92.0000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 53.8500 91.4000 53.9500 92.0000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 52.2500 91.4000 52.3500 92.0000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 50.6500 91.4000 50.7500 92.0000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 49.0500 91.4000 49.1500 92.0000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 47.4500 91.4000 47.5500 92.0000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 45.8500 91.4000 45.9500 92.0000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 44.2500 91.4000 44.3500 92.0000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 42.6500 91.4000 42.7500 92.0000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 41.0500 91.4000 41.1500 92.0000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 39.4500 91.4000 39.5500 92.0000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 37.8500 91.4000 37.9500 92.0000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 36.2500 91.4000 36.3500 92.0000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 34.6500 91.4000 34.7500 92.0000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 33.0500 91.4000 33.1500 92.0000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 31.4500 91.4000 31.5500 92.0000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 29.8500 91.4000 29.9500 92.0000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 28.2500 91.4000 28.3500 92.0000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 26.6500 91.4000 26.7500 92.0000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 25.0500 91.4000 25.1500 92.0000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 42.1500 0.6000 42.2500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.1500 0.6000 34.2500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 46.1500 0.6000 46.2500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 50.1500 0.6000 50.2500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 54.1500 0.6000 54.2500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 58.1500 0.6000 58.2500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 228.9900 10.0000 230.9900 82.0000 ;
        RECT 162.6600 10.0000 164.6600 82.0000 ;
        RECT 96.3300 10.0000 98.3300 82.0000 ;
        RECT 30.0000 10.0000 32.0000 82.0000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 235.9900 10.0000 237.9900 82.0000 ;
        RECT 169.6600 10.0000 171.6600 82.0000 ;
        RECT 103.3300 10.0000 105.3300 82.0000 ;
        RECT 37.0000 10.0000 39.0000 82.0000 ;
        RECT 37.0000 9.8350 39.0000 10.1650 ;
        RECT 103.3300 9.8350 105.3300 10.1650 ;
        RECT 169.6600 9.8350 171.6600 10.1650 ;
        RECT 235.9900 9.8350 237.9900 10.1650 ;
        RECT 37.0000 81.8350 39.0000 82.1650 ;
        RECT 103.3300 81.8350 105.3300 82.1650 ;
        RECT 169.6600 81.8350 171.6600 82.1650 ;
        RECT 235.9900 81.8350 237.9900 82.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 268.0000 92.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 268.0000 92.0000 ;
    LAYER M3 ;
      RECT 228.5100 91.2400 268.0000 92.0000 ;
      RECT 226.9100 91.2400 228.0900 92.0000 ;
      RECT 225.3100 91.2400 226.4900 92.0000 ;
      RECT 223.7100 91.2400 224.8900 92.0000 ;
      RECT 222.1100 91.2400 223.2900 92.0000 ;
      RECT 220.5100 91.2400 221.6900 92.0000 ;
      RECT 218.9100 91.2400 220.0900 92.0000 ;
      RECT 217.3100 91.2400 218.4900 92.0000 ;
      RECT 215.7100 91.2400 216.8900 92.0000 ;
      RECT 214.1100 91.2400 215.2900 92.0000 ;
      RECT 212.5100 91.2400 213.6900 92.0000 ;
      RECT 210.9100 91.2400 212.0900 92.0000 ;
      RECT 209.3100 91.2400 210.4900 92.0000 ;
      RECT 207.7100 91.2400 208.8900 92.0000 ;
      RECT 206.1100 91.2400 207.2900 92.0000 ;
      RECT 204.5100 91.2400 205.6900 92.0000 ;
      RECT 202.9100 91.2400 204.0900 92.0000 ;
      RECT 201.3100 91.2400 202.4900 92.0000 ;
      RECT 199.7100 91.2400 200.8900 92.0000 ;
      RECT 198.1100 91.2400 199.2900 92.0000 ;
      RECT 196.5100 91.2400 197.6900 92.0000 ;
      RECT 194.9100 91.2400 196.0900 92.0000 ;
      RECT 193.3100 91.2400 194.4900 92.0000 ;
      RECT 191.7100 91.2400 192.8900 92.0000 ;
      RECT 190.1100 91.2400 191.2900 92.0000 ;
      RECT 188.5100 91.2400 189.6900 92.0000 ;
      RECT 186.9100 91.2400 188.0900 92.0000 ;
      RECT 185.3100 91.2400 186.4900 92.0000 ;
      RECT 183.7100 91.2400 184.8900 92.0000 ;
      RECT 182.1100 91.2400 183.2900 92.0000 ;
      RECT 180.5100 91.2400 181.6900 92.0000 ;
      RECT 178.9100 91.2400 180.0900 92.0000 ;
      RECT 177.3100 91.2400 178.4900 92.0000 ;
      RECT 175.7100 91.2400 176.8900 92.0000 ;
      RECT 174.1100 91.2400 175.2900 92.0000 ;
      RECT 172.5100 91.2400 173.6900 92.0000 ;
      RECT 170.9100 91.2400 172.0900 92.0000 ;
      RECT 169.3100 91.2400 170.4900 92.0000 ;
      RECT 167.7100 91.2400 168.8900 92.0000 ;
      RECT 166.1100 91.2400 167.2900 92.0000 ;
      RECT 164.5100 91.2400 165.6900 92.0000 ;
      RECT 162.9100 91.2400 164.0900 92.0000 ;
      RECT 161.3100 91.2400 162.4900 92.0000 ;
      RECT 159.7100 91.2400 160.8900 92.0000 ;
      RECT 158.1100 91.2400 159.2900 92.0000 ;
      RECT 156.5100 91.2400 157.6900 92.0000 ;
      RECT 154.9100 91.2400 156.0900 92.0000 ;
      RECT 153.3100 91.2400 154.4900 92.0000 ;
      RECT 151.7100 91.2400 152.8900 92.0000 ;
      RECT 150.1100 91.2400 151.2900 92.0000 ;
      RECT 148.5100 91.2400 149.6900 92.0000 ;
      RECT 146.9100 91.2400 148.0900 92.0000 ;
      RECT 145.3100 91.2400 146.4900 92.0000 ;
      RECT 143.7100 91.2400 144.8900 92.0000 ;
      RECT 142.1100 91.2400 143.2900 92.0000 ;
      RECT 140.5100 91.2400 141.6900 92.0000 ;
      RECT 138.9100 91.2400 140.0900 92.0000 ;
      RECT 137.3100 91.2400 138.4900 92.0000 ;
      RECT 135.7100 91.2400 136.8900 92.0000 ;
      RECT 134.1100 91.2400 135.2900 92.0000 ;
      RECT 132.5100 91.2400 133.6900 92.0000 ;
      RECT 130.9100 91.2400 132.0900 92.0000 ;
      RECT 129.3100 91.2400 130.4900 92.0000 ;
      RECT 127.7100 91.2400 128.8900 92.0000 ;
      RECT 126.1100 91.2400 127.2900 92.0000 ;
      RECT 124.5100 91.2400 125.6900 92.0000 ;
      RECT 122.9100 91.2400 124.0900 92.0000 ;
      RECT 121.3100 91.2400 122.4900 92.0000 ;
      RECT 119.7100 91.2400 120.8900 92.0000 ;
      RECT 118.1100 91.2400 119.2900 92.0000 ;
      RECT 116.5100 91.2400 117.6900 92.0000 ;
      RECT 114.9100 91.2400 116.0900 92.0000 ;
      RECT 113.3100 91.2400 114.4900 92.0000 ;
      RECT 111.7100 91.2400 112.8900 92.0000 ;
      RECT 110.1100 91.2400 111.2900 92.0000 ;
      RECT 108.5100 91.2400 109.6900 92.0000 ;
      RECT 106.9100 91.2400 108.0900 92.0000 ;
      RECT 105.3100 91.2400 106.4900 92.0000 ;
      RECT 103.7100 91.2400 104.8900 92.0000 ;
      RECT 102.1100 91.2400 103.2900 92.0000 ;
      RECT 100.5100 91.2400 101.6900 92.0000 ;
      RECT 98.9100 91.2400 100.0900 92.0000 ;
      RECT 97.3100 91.2400 98.4900 92.0000 ;
      RECT 95.7100 91.2400 96.8900 92.0000 ;
      RECT 94.1100 91.2400 95.2900 92.0000 ;
      RECT 92.5100 91.2400 93.6900 92.0000 ;
      RECT 90.9100 91.2400 92.0900 92.0000 ;
      RECT 89.3100 91.2400 90.4900 92.0000 ;
      RECT 87.7100 91.2400 88.8900 92.0000 ;
      RECT 86.1100 91.2400 87.2900 92.0000 ;
      RECT 84.5100 91.2400 85.6900 92.0000 ;
      RECT 82.9100 91.2400 84.0900 92.0000 ;
      RECT 81.3100 91.2400 82.4900 92.0000 ;
      RECT 79.7100 91.2400 80.8900 92.0000 ;
      RECT 78.1100 91.2400 79.2900 92.0000 ;
      RECT 76.5100 91.2400 77.6900 92.0000 ;
      RECT 74.9100 91.2400 76.0900 92.0000 ;
      RECT 73.3100 91.2400 74.4900 92.0000 ;
      RECT 71.7100 91.2400 72.8900 92.0000 ;
      RECT 70.1100 91.2400 71.2900 92.0000 ;
      RECT 68.5100 91.2400 69.6900 92.0000 ;
      RECT 66.9100 91.2400 68.0900 92.0000 ;
      RECT 65.3100 91.2400 66.4900 92.0000 ;
      RECT 63.7100 91.2400 64.8900 92.0000 ;
      RECT 62.1100 91.2400 63.2900 92.0000 ;
      RECT 60.5100 91.2400 61.6900 92.0000 ;
      RECT 58.9100 91.2400 60.0900 92.0000 ;
      RECT 57.3100 91.2400 58.4900 92.0000 ;
      RECT 55.7100 91.2400 56.8900 92.0000 ;
      RECT 54.1100 91.2400 55.2900 92.0000 ;
      RECT 52.5100 91.2400 53.6900 92.0000 ;
      RECT 50.9100 91.2400 52.0900 92.0000 ;
      RECT 49.3100 91.2400 50.4900 92.0000 ;
      RECT 47.7100 91.2400 48.8900 92.0000 ;
      RECT 46.1100 91.2400 47.2900 92.0000 ;
      RECT 44.5100 91.2400 45.6900 92.0000 ;
      RECT 42.9100 91.2400 44.0900 92.0000 ;
      RECT 41.3100 91.2400 42.4900 92.0000 ;
      RECT 39.7100 91.2400 40.8900 92.0000 ;
      RECT 38.1100 91.2400 39.2900 92.0000 ;
      RECT 36.5100 91.2400 37.6900 92.0000 ;
      RECT 34.9100 91.2400 36.0900 92.0000 ;
      RECT 33.3100 91.2400 34.4900 92.0000 ;
      RECT 31.7100 91.2400 32.8900 92.0000 ;
      RECT 30.1100 91.2400 31.2900 92.0000 ;
      RECT 28.5100 91.2400 29.6900 92.0000 ;
      RECT 26.9100 91.2400 28.0900 92.0000 ;
      RECT 25.3100 91.2400 26.4900 92.0000 ;
      RECT 0.0000 91.2400 24.8900 92.0000 ;
      RECT 0.0000 58.3500 268.0000 91.2400 ;
      RECT 0.7000 58.0500 268.0000 58.3500 ;
      RECT 0.0000 54.3500 268.0000 58.0500 ;
      RECT 0.7000 54.0500 268.0000 54.3500 ;
      RECT 0.0000 50.3500 268.0000 54.0500 ;
      RECT 0.7000 50.0500 268.0000 50.3500 ;
      RECT 0.0000 46.3500 268.0000 50.0500 ;
      RECT 0.7000 46.0500 268.0000 46.3500 ;
      RECT 0.0000 42.3500 268.0000 46.0500 ;
      RECT 0.7000 42.0500 268.0000 42.3500 ;
      RECT 0.0000 38.3500 268.0000 42.0500 ;
      RECT 0.7000 38.0500 268.0000 38.3500 ;
      RECT 0.0000 34.3500 268.0000 38.0500 ;
      RECT 0.7000 34.0500 268.0000 34.3500 ;
      RECT 0.0000 0.7600 268.0000 34.0500 ;
      RECT 228.5100 0.0000 268.0000 0.7600 ;
      RECT 226.9100 0.0000 228.0900 0.7600 ;
      RECT 225.3100 0.0000 226.4900 0.7600 ;
      RECT 223.7100 0.0000 224.8900 0.7600 ;
      RECT 222.1100 0.0000 223.2900 0.7600 ;
      RECT 220.5100 0.0000 221.6900 0.7600 ;
      RECT 218.9100 0.0000 220.0900 0.7600 ;
      RECT 217.3100 0.0000 218.4900 0.7600 ;
      RECT 215.7100 0.0000 216.8900 0.7600 ;
      RECT 214.1100 0.0000 215.2900 0.7600 ;
      RECT 212.5100 0.0000 213.6900 0.7600 ;
      RECT 210.9100 0.0000 212.0900 0.7600 ;
      RECT 209.3100 0.0000 210.4900 0.7600 ;
      RECT 207.7100 0.0000 208.8900 0.7600 ;
      RECT 206.1100 0.0000 207.2900 0.7600 ;
      RECT 204.5100 0.0000 205.6900 0.7600 ;
      RECT 202.9100 0.0000 204.0900 0.7600 ;
      RECT 201.3100 0.0000 202.4900 0.7600 ;
      RECT 199.7100 0.0000 200.8900 0.7600 ;
      RECT 198.1100 0.0000 199.2900 0.7600 ;
      RECT 196.5100 0.0000 197.6900 0.7600 ;
      RECT 194.9100 0.0000 196.0900 0.7600 ;
      RECT 193.3100 0.0000 194.4900 0.7600 ;
      RECT 191.7100 0.0000 192.8900 0.7600 ;
      RECT 190.1100 0.0000 191.2900 0.7600 ;
      RECT 188.5100 0.0000 189.6900 0.7600 ;
      RECT 186.9100 0.0000 188.0900 0.7600 ;
      RECT 185.3100 0.0000 186.4900 0.7600 ;
      RECT 183.7100 0.0000 184.8900 0.7600 ;
      RECT 182.1100 0.0000 183.2900 0.7600 ;
      RECT 180.5100 0.0000 181.6900 0.7600 ;
      RECT 178.9100 0.0000 180.0900 0.7600 ;
      RECT 177.3100 0.0000 178.4900 0.7600 ;
      RECT 175.7100 0.0000 176.8900 0.7600 ;
      RECT 174.1100 0.0000 175.2900 0.7600 ;
      RECT 172.5100 0.0000 173.6900 0.7600 ;
      RECT 170.9100 0.0000 172.0900 0.7600 ;
      RECT 169.3100 0.0000 170.4900 0.7600 ;
      RECT 167.7100 0.0000 168.8900 0.7600 ;
      RECT 166.1100 0.0000 167.2900 0.7600 ;
      RECT 164.5100 0.0000 165.6900 0.7600 ;
      RECT 162.9100 0.0000 164.0900 0.7600 ;
      RECT 161.3100 0.0000 162.4900 0.7600 ;
      RECT 159.7100 0.0000 160.8900 0.7600 ;
      RECT 158.1100 0.0000 159.2900 0.7600 ;
      RECT 156.5100 0.0000 157.6900 0.7600 ;
      RECT 154.9100 0.0000 156.0900 0.7600 ;
      RECT 153.3100 0.0000 154.4900 0.7600 ;
      RECT 151.7100 0.0000 152.8900 0.7600 ;
      RECT 150.1100 0.0000 151.2900 0.7600 ;
      RECT 148.5100 0.0000 149.6900 0.7600 ;
      RECT 146.9100 0.0000 148.0900 0.7600 ;
      RECT 145.3100 0.0000 146.4900 0.7600 ;
      RECT 143.7100 0.0000 144.8900 0.7600 ;
      RECT 142.1100 0.0000 143.2900 0.7600 ;
      RECT 140.5100 0.0000 141.6900 0.7600 ;
      RECT 138.9100 0.0000 140.0900 0.7600 ;
      RECT 137.3100 0.0000 138.4900 0.7600 ;
      RECT 135.7100 0.0000 136.8900 0.7600 ;
      RECT 134.1100 0.0000 135.2900 0.7600 ;
      RECT 132.5100 0.0000 133.6900 0.7600 ;
      RECT 130.9100 0.0000 132.0900 0.7600 ;
      RECT 129.3100 0.0000 130.4900 0.7600 ;
      RECT 127.7100 0.0000 128.8900 0.7600 ;
      RECT 126.1100 0.0000 127.2900 0.7600 ;
      RECT 124.5100 0.0000 125.6900 0.7600 ;
      RECT 122.9100 0.0000 124.0900 0.7600 ;
      RECT 121.3100 0.0000 122.4900 0.7600 ;
      RECT 119.7100 0.0000 120.8900 0.7600 ;
      RECT 118.1100 0.0000 119.2900 0.7600 ;
      RECT 116.5100 0.0000 117.6900 0.7600 ;
      RECT 114.9100 0.0000 116.0900 0.7600 ;
      RECT 113.3100 0.0000 114.4900 0.7600 ;
      RECT 111.7100 0.0000 112.8900 0.7600 ;
      RECT 110.1100 0.0000 111.2900 0.7600 ;
      RECT 108.5100 0.0000 109.6900 0.7600 ;
      RECT 106.9100 0.0000 108.0900 0.7600 ;
      RECT 105.3100 0.0000 106.4900 0.7600 ;
      RECT 103.7100 0.0000 104.8900 0.7600 ;
      RECT 102.1100 0.0000 103.2900 0.7600 ;
      RECT 100.5100 0.0000 101.6900 0.7600 ;
      RECT 98.9100 0.0000 100.0900 0.7600 ;
      RECT 97.3100 0.0000 98.4900 0.7600 ;
      RECT 95.7100 0.0000 96.8900 0.7600 ;
      RECT 94.1100 0.0000 95.2900 0.7600 ;
      RECT 92.5100 0.0000 93.6900 0.7600 ;
      RECT 90.9100 0.0000 92.0900 0.7600 ;
      RECT 89.3100 0.0000 90.4900 0.7600 ;
      RECT 87.7100 0.0000 88.8900 0.7600 ;
      RECT 86.1100 0.0000 87.2900 0.7600 ;
      RECT 84.5100 0.0000 85.6900 0.7600 ;
      RECT 82.9100 0.0000 84.0900 0.7600 ;
      RECT 81.3100 0.0000 82.4900 0.7600 ;
      RECT 79.7100 0.0000 80.8900 0.7600 ;
      RECT 78.1100 0.0000 79.2900 0.7600 ;
      RECT 76.5100 0.0000 77.6900 0.7600 ;
      RECT 74.9100 0.0000 76.0900 0.7600 ;
      RECT 73.3100 0.0000 74.4900 0.7600 ;
      RECT 71.7100 0.0000 72.8900 0.7600 ;
      RECT 70.1100 0.0000 71.2900 0.7600 ;
      RECT 68.5100 0.0000 69.6900 0.7600 ;
      RECT 66.9100 0.0000 68.0900 0.7600 ;
      RECT 65.3100 0.0000 66.4900 0.7600 ;
      RECT 63.7100 0.0000 64.8900 0.7600 ;
      RECT 62.1100 0.0000 63.2900 0.7600 ;
      RECT 60.5100 0.0000 61.6900 0.7600 ;
      RECT 58.9100 0.0000 60.0900 0.7600 ;
      RECT 57.3100 0.0000 58.4900 0.7600 ;
      RECT 55.7100 0.0000 56.8900 0.7600 ;
      RECT 54.1100 0.0000 55.2900 0.7600 ;
      RECT 52.5100 0.0000 53.6900 0.7600 ;
      RECT 50.9100 0.0000 52.0900 0.7600 ;
      RECT 49.3100 0.0000 50.4900 0.7600 ;
      RECT 47.7100 0.0000 48.8900 0.7600 ;
      RECT 46.1100 0.0000 47.2900 0.7600 ;
      RECT 44.5100 0.0000 45.6900 0.7600 ;
      RECT 42.9100 0.0000 44.0900 0.7600 ;
      RECT 41.3100 0.0000 42.4900 0.7600 ;
      RECT 39.7100 0.0000 40.8900 0.7600 ;
      RECT 38.1100 0.0000 39.2900 0.7600 ;
      RECT 36.5100 0.0000 37.6900 0.7600 ;
      RECT 34.9100 0.0000 36.0900 0.7600 ;
      RECT 33.3100 0.0000 34.4900 0.7600 ;
      RECT 31.7100 0.0000 32.8900 0.7600 ;
      RECT 30.1100 0.0000 31.2900 0.7600 ;
      RECT 28.5100 0.0000 29.6900 0.7600 ;
      RECT 26.9100 0.0000 28.0900 0.7600 ;
      RECT 25.3100 0.0000 26.4900 0.7600 ;
      RECT 0.0000 0.0000 24.8900 0.7600 ;
    LAYER M4 ;
      RECT 0.0000 82.6650 268.0000 92.0000 ;
      RECT 172.1600 82.5000 235.4900 82.6650 ;
      RECT 105.8300 82.5000 169.1600 82.6650 ;
      RECT 39.5000 82.5000 102.8300 82.6650 ;
      RECT 0.0000 82.5000 36.5000 82.6650 ;
      RECT 231.4900 9.5000 235.4900 82.5000 ;
      RECT 172.1600 9.5000 228.4900 82.5000 ;
      RECT 165.1600 9.5000 169.1600 82.5000 ;
      RECT 105.8300 9.5000 162.1600 82.5000 ;
      RECT 98.8300 9.5000 102.8300 82.5000 ;
      RECT 39.5000 9.5000 95.8300 82.5000 ;
      RECT 32.5000 9.5000 36.5000 82.5000 ;
      RECT 0.0000 9.5000 29.5000 82.5000 ;
      RECT 238.4900 9.3350 268.0000 82.6650 ;
      RECT 172.1600 9.3350 235.4900 9.5000 ;
      RECT 105.8300 9.3350 169.1600 9.5000 ;
      RECT 39.5000 9.3350 102.8300 9.5000 ;
      RECT 0.0000 9.3350 36.5000 9.5000 ;
      RECT 0.0000 0.0000 268.0000 9.3350 ;
  END
END sram_w16

END LIBRARY
