##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 22 18:56:50 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 608.8000 BY 311.6000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 81.7500 0.5200 81.8500 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 227.5500 0.5200 227.6500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 225.7500 0.5200 225.8500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 223.9500 0.5200 224.0500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 222.1500 0.5200 222.2500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 220.3500 0.5200 220.4500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 218.5500 0.5200 218.6500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 216.7500 0.5200 216.8500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 214.9500 0.5200 215.0500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 213.1500 0.5200 213.2500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 211.3500 0.5200 211.4500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 209.5500 0.5200 209.6500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 207.7500 0.5200 207.8500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 205.9500 0.5200 206.0500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 204.1500 0.5200 204.2500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 202.3500 0.5200 202.4500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 200.5500 0.5200 200.6500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 198.7500 0.5200 198.8500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 196.9500 0.5200 197.0500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 195.1500 0.5200 195.2500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 193.3500 0.5200 193.4500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 191.5500 0.5200 191.6500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 189.7500 0.5200 189.8500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 187.9500 0.5200 188.0500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 186.1500 0.5200 186.2500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 184.3500 0.5200 184.4500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 182.5500 0.5200 182.6500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 180.7500 0.5200 180.8500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 178.9500 0.5200 179.0500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 177.1500 0.5200 177.2500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 175.3500 0.5200 175.4500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 173.5500 0.5200 173.6500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 171.7500 0.5200 171.8500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 169.9500 0.5200 170.0500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 168.1500 0.5200 168.2500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 166.3500 0.5200 166.4500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 164.5500 0.5200 164.6500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 162.7500 0.5200 162.8500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 160.9500 0.5200 161.0500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 159.1500 0.5200 159.2500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 157.3500 0.5200 157.4500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 155.5500 0.5200 155.6500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 153.7500 0.5200 153.8500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 151.9500 0.5200 152.0500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 150.1500 0.5200 150.2500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 148.3500 0.5200 148.4500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 146.5500 0.5200 146.6500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 144.7500 0.5200 144.8500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 142.9500 0.5200 143.0500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 141.1500 0.5200 141.2500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 139.3500 0.5200 139.4500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 137.5500 0.5200 137.6500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 135.7500 0.5200 135.8500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 133.9500 0.5200 134.0500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 132.1500 0.5200 132.2500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 130.3500 0.5200 130.4500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 128.5500 0.5200 128.6500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 126.7500 0.5200 126.8500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 124.9500 0.5200 125.0500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 123.1500 0.5200 123.2500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 121.3500 0.5200 121.4500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 119.5500 0.5200 119.6500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 117.7500 0.5200 117.8500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 115.9500 0.5200 116.0500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 114.1500 0.5200 114.2500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.2500 0.0000 18.3500 0.5200 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.8500 0.0000 21.9500 0.5200 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.4500 0.0000 25.5500 0.5200 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.0500 0.0000 29.1500 0.5200 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.6500 0.0000 32.7500 0.5200 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.2500 0.0000 36.3500 0.5200 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.8500 0.0000 39.9500 0.5200 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.4500 0.0000 43.5500 0.5200 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.0500 0.0000 47.1500 0.5200 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.6500 0.0000 50.7500 0.5200 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.2500 0.0000 54.3500 0.5200 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.8500 0.0000 57.9500 0.5200 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.4500 0.0000 61.5500 0.5200 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.0500 0.0000 65.1500 0.5200 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.6500 0.0000 68.7500 0.5200 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.2500 0.0000 72.3500 0.5200 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.8500 0.0000 75.9500 0.5200 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.4500 0.0000 79.5500 0.5200 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.0500 0.0000 83.1500 0.5200 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.6500 0.0000 86.7500 0.5200 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.2500 0.0000 90.3500 0.5200 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.8500 0.0000 93.9500 0.5200 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.4500 0.0000 97.5500 0.5200 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.0500 0.0000 101.1500 0.5200 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.6500 0.0000 104.7500 0.5200 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.2500 0.0000 108.3500 0.5200 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.8500 0.0000 111.9500 0.5200 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.4500 0.0000 115.5500 0.5200 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.0500 0.0000 119.1500 0.5200 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.6500 0.0000 122.7500 0.5200 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.2500 0.0000 126.3500 0.5200 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.8500 0.0000 129.9500 0.5200 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.4500 0.0000 133.5500 0.5200 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.0500 0.0000 137.1500 0.5200 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.6500 0.0000 140.7500 0.5200 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.2500 0.0000 144.3500 0.5200 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.8500 0.0000 147.9500 0.5200 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.4500 0.0000 151.5500 0.5200 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.0500 0.0000 155.1500 0.5200 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.6500 0.0000 158.7500 0.5200 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.2500 0.0000 162.3500 0.5200 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.8500 0.0000 165.9500 0.5200 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.4500 0.0000 169.5500 0.5200 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.0500 0.0000 173.1500 0.5200 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.6500 0.0000 176.7500 0.5200 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.2500 0.0000 180.3500 0.5200 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.8500 0.0000 183.9500 0.5200 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.4500 0.0000 187.5500 0.5200 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.0500 0.0000 191.1500 0.5200 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.6500 0.0000 194.7500 0.5200 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.2500 0.0000 198.3500 0.5200 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.8500 0.0000 201.9500 0.5200 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.4500 0.0000 205.5500 0.5200 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.0500 0.0000 209.1500 0.5200 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.6500 0.0000 212.7500 0.5200 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.2500 0.0000 216.3500 0.5200 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.8500 0.0000 219.9500 0.5200 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.4500 0.0000 223.5500 0.5200 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.0500 0.0000 227.1500 0.5200 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.6500 0.0000 230.7500 0.5200 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.2500 0.0000 234.3500 0.5200 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.8500 0.0000 237.9500 0.5200 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.4500 0.0000 241.5500 0.5200 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 245.0500 0.0000 245.1500 0.5200 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.6500 0.0000 248.7500 0.5200 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.2500 0.0000 252.3500 0.5200 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.8500 0.0000 255.9500 0.5200 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.4500 0.0000 259.5500 0.5200 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.0500 0.0000 263.1500 0.5200 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 266.6500 0.0000 266.7500 0.5200 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.2500 0.0000 270.3500 0.5200 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.8500 0.0000 273.9500 0.5200 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.4500 0.0000 277.5500 0.5200 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.0500 0.0000 281.1500 0.5200 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284.6500 0.0000 284.7500 0.5200 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.2500 0.0000 288.3500 0.5200 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.8500 0.0000 291.9500 0.5200 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.4500 0.0000 295.5500 0.5200 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.0500 0.0000 299.1500 0.5200 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.6500 0.0000 302.7500 0.5200 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.2500 0.0000 306.3500 0.5200 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.8500 0.0000 309.9500 0.5200 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.4500 0.0000 313.5500 0.5200 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.0500 0.0000 317.1500 0.5200 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.6500 0.0000 320.7500 0.5200 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.2500 0.0000 324.3500 0.5200 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.8500 0.0000 327.9500 0.5200 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.4500 0.0000 331.5500 0.5200 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.0500 0.0000 335.1500 0.5200 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.6500 0.0000 338.7500 0.5200 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.2500 0.0000 342.3500 0.5200 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.8500 0.0000 345.9500 0.5200 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.4500 0.0000 349.5500 0.5200 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.0500 0.0000 353.1500 0.5200 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.6500 0.0000 356.7500 0.5200 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.2500 0.0000 360.3500 0.5200 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.8500 0.0000 363.9500 0.5200 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.4500 0.0000 367.5500 0.5200 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.0500 0.0000 371.1500 0.5200 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.6500 0.0000 374.7500 0.5200 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.2500 0.0000 378.3500 0.5200 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.8500 0.0000 381.9500 0.5200 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 385.4500 0.0000 385.5500 0.5200 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 389.0500 0.0000 389.1500 0.5200 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.6500 0.0000 392.7500 0.5200 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.2500 0.0000 396.3500 0.5200 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.8500 0.0000 399.9500 0.5200 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.4500 0.0000 403.5500 0.5200 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.0500 0.0000 407.1500 0.5200 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.6500 0.0000 410.7500 0.5200 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.2500 0.0000 414.3500 0.5200 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.8500 0.0000 417.9500 0.5200 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 421.4500 0.0000 421.5500 0.5200 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 425.0500 0.0000 425.1500 0.5200 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.6500 0.0000 428.7500 0.5200 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.2500 0.0000 432.3500 0.5200 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.8500 0.0000 435.9500 0.5200 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.4500 0.0000 439.5500 0.5200 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.0500 0.0000 443.1500 0.5200 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 446.6500 0.0000 446.7500 0.5200 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.2500 0.0000 450.3500 0.5200 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 453.8500 0.0000 453.9500 0.5200 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.4500 0.0000 457.5500 0.5200 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 461.0500 0.0000 461.1500 0.5200 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 464.6500 0.0000 464.7500 0.5200 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 468.2500 0.0000 468.3500 0.5200 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 471.8500 0.0000 471.9500 0.5200 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 475.4500 0.0000 475.5500 0.5200 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 479.0500 0.0000 479.1500 0.5200 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 482.6500 0.0000 482.7500 0.5200 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 486.2500 0.0000 486.3500 0.5200 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 489.8500 0.0000 489.9500 0.5200 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 493.4500 0.0000 493.5500 0.5200 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 497.0500 0.0000 497.1500 0.5200 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 500.6500 0.0000 500.7500 0.5200 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 504.2500 0.0000 504.3500 0.5200 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 507.8500 0.0000 507.9500 0.5200 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 511.4500 0.0000 511.5500 0.5200 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 515.0500 0.0000 515.1500 0.5200 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 518.6500 0.0000 518.7500 0.5200 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 522.2500 0.0000 522.3500 0.5200 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 525.8500 0.0000 525.9500 0.5200 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 529.4500 0.0000 529.5500 0.5200 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 533.0500 0.0000 533.1500 0.5200 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.6500 0.0000 536.7500 0.5200 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 540.2500 0.0000 540.3500 0.5200 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 543.8500 0.0000 543.9500 0.5200 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 547.4500 0.0000 547.5500 0.5200 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 551.0500 0.0000 551.1500 0.5200 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 554.6500 0.0000 554.7500 0.5200 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 558.2500 0.0000 558.3500 0.5200 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 561.8500 0.0000 561.9500 0.5200 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 565.4500 0.0000 565.5500 0.5200 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 569.0500 0.0000 569.1500 0.5200 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 572.6500 0.0000 572.7500 0.5200 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 576.2500 0.0000 576.3500 0.5200 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 579.8500 0.0000 579.9500 0.5200 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 583.4500 0.0000 583.5500 0.5200 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 587.0500 0.0000 587.1500 0.5200 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 590.6500 0.0000 590.7500 0.5200 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 112.3500 0.5200 112.4500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 110.5500 0.5200 110.6500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 108.7500 0.5200 108.8500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 106.9500 0.5200 107.0500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 105.1500 0.5200 105.2500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 103.3500 0.5200 103.4500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 101.5500 0.5200 101.6500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 99.7500 0.5200 99.8500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 97.9500 0.5200 98.0500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 96.1500 0.5200 96.2500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 94.3500 0.5200 94.4500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 92.5500 0.5200 92.6500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 90.7500 0.5200 90.8500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 88.9500 0.5200 89.0500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 87.1500 0.5200 87.2500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 85.3500 0.5200 85.4500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 83.5500 0.5200 83.6500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 229.3500 0.5200 229.4500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 608.8000 311.6000 ;
    LAYER M2 ;
      RECT 0.0000 0.6200 608.8000 311.6000 ;
      RECT 590.8500 0.0000 608.8000 0.6200 ;
      RECT 587.2500 0.0000 590.5500 0.6200 ;
      RECT 583.6500 0.0000 586.9500 0.6200 ;
      RECT 580.0500 0.0000 583.3500 0.6200 ;
      RECT 576.4500 0.0000 579.7500 0.6200 ;
      RECT 572.8500 0.0000 576.1500 0.6200 ;
      RECT 569.2500 0.0000 572.5500 0.6200 ;
      RECT 565.6500 0.0000 568.9500 0.6200 ;
      RECT 562.0500 0.0000 565.3500 0.6200 ;
      RECT 558.4500 0.0000 561.7500 0.6200 ;
      RECT 554.8500 0.0000 558.1500 0.6200 ;
      RECT 551.2500 0.0000 554.5500 0.6200 ;
      RECT 547.6500 0.0000 550.9500 0.6200 ;
      RECT 544.0500 0.0000 547.3500 0.6200 ;
      RECT 540.4500 0.0000 543.7500 0.6200 ;
      RECT 536.8500 0.0000 540.1500 0.6200 ;
      RECT 533.2500 0.0000 536.5500 0.6200 ;
      RECT 529.6500 0.0000 532.9500 0.6200 ;
      RECT 526.0500 0.0000 529.3500 0.6200 ;
      RECT 522.4500 0.0000 525.7500 0.6200 ;
      RECT 518.8500 0.0000 522.1500 0.6200 ;
      RECT 515.2500 0.0000 518.5500 0.6200 ;
      RECT 511.6500 0.0000 514.9500 0.6200 ;
      RECT 508.0500 0.0000 511.3500 0.6200 ;
      RECT 504.4500 0.0000 507.7500 0.6200 ;
      RECT 500.8500 0.0000 504.1500 0.6200 ;
      RECT 497.2500 0.0000 500.5500 0.6200 ;
      RECT 493.6500 0.0000 496.9500 0.6200 ;
      RECT 490.0500 0.0000 493.3500 0.6200 ;
      RECT 486.4500 0.0000 489.7500 0.6200 ;
      RECT 482.8500 0.0000 486.1500 0.6200 ;
      RECT 479.2500 0.0000 482.5500 0.6200 ;
      RECT 475.6500 0.0000 478.9500 0.6200 ;
      RECT 472.0500 0.0000 475.3500 0.6200 ;
      RECT 468.4500 0.0000 471.7500 0.6200 ;
      RECT 464.8500 0.0000 468.1500 0.6200 ;
      RECT 461.2500 0.0000 464.5500 0.6200 ;
      RECT 457.6500 0.0000 460.9500 0.6200 ;
      RECT 454.0500 0.0000 457.3500 0.6200 ;
      RECT 450.4500 0.0000 453.7500 0.6200 ;
      RECT 446.8500 0.0000 450.1500 0.6200 ;
      RECT 443.2500 0.0000 446.5500 0.6200 ;
      RECT 439.6500 0.0000 442.9500 0.6200 ;
      RECT 436.0500 0.0000 439.3500 0.6200 ;
      RECT 432.4500 0.0000 435.7500 0.6200 ;
      RECT 428.8500 0.0000 432.1500 0.6200 ;
      RECT 425.2500 0.0000 428.5500 0.6200 ;
      RECT 421.6500 0.0000 424.9500 0.6200 ;
      RECT 418.0500 0.0000 421.3500 0.6200 ;
      RECT 414.4500 0.0000 417.7500 0.6200 ;
      RECT 410.8500 0.0000 414.1500 0.6200 ;
      RECT 407.2500 0.0000 410.5500 0.6200 ;
      RECT 403.6500 0.0000 406.9500 0.6200 ;
      RECT 400.0500 0.0000 403.3500 0.6200 ;
      RECT 396.4500 0.0000 399.7500 0.6200 ;
      RECT 392.8500 0.0000 396.1500 0.6200 ;
      RECT 389.2500 0.0000 392.5500 0.6200 ;
      RECT 385.6500 0.0000 388.9500 0.6200 ;
      RECT 382.0500 0.0000 385.3500 0.6200 ;
      RECT 378.4500 0.0000 381.7500 0.6200 ;
      RECT 374.8500 0.0000 378.1500 0.6200 ;
      RECT 371.2500 0.0000 374.5500 0.6200 ;
      RECT 367.6500 0.0000 370.9500 0.6200 ;
      RECT 364.0500 0.0000 367.3500 0.6200 ;
      RECT 360.4500 0.0000 363.7500 0.6200 ;
      RECT 356.8500 0.0000 360.1500 0.6200 ;
      RECT 353.2500 0.0000 356.5500 0.6200 ;
      RECT 349.6500 0.0000 352.9500 0.6200 ;
      RECT 346.0500 0.0000 349.3500 0.6200 ;
      RECT 342.4500 0.0000 345.7500 0.6200 ;
      RECT 338.8500 0.0000 342.1500 0.6200 ;
      RECT 335.2500 0.0000 338.5500 0.6200 ;
      RECT 331.6500 0.0000 334.9500 0.6200 ;
      RECT 328.0500 0.0000 331.3500 0.6200 ;
      RECT 324.4500 0.0000 327.7500 0.6200 ;
      RECT 320.8500 0.0000 324.1500 0.6200 ;
      RECT 317.2500 0.0000 320.5500 0.6200 ;
      RECT 313.6500 0.0000 316.9500 0.6200 ;
      RECT 310.0500 0.0000 313.3500 0.6200 ;
      RECT 306.4500 0.0000 309.7500 0.6200 ;
      RECT 302.8500 0.0000 306.1500 0.6200 ;
      RECT 299.2500 0.0000 302.5500 0.6200 ;
      RECT 295.6500 0.0000 298.9500 0.6200 ;
      RECT 292.0500 0.0000 295.3500 0.6200 ;
      RECT 288.4500 0.0000 291.7500 0.6200 ;
      RECT 284.8500 0.0000 288.1500 0.6200 ;
      RECT 281.2500 0.0000 284.5500 0.6200 ;
      RECT 277.6500 0.0000 280.9500 0.6200 ;
      RECT 274.0500 0.0000 277.3500 0.6200 ;
      RECT 270.4500 0.0000 273.7500 0.6200 ;
      RECT 266.8500 0.0000 270.1500 0.6200 ;
      RECT 263.2500 0.0000 266.5500 0.6200 ;
      RECT 259.6500 0.0000 262.9500 0.6200 ;
      RECT 256.0500 0.0000 259.3500 0.6200 ;
      RECT 252.4500 0.0000 255.7500 0.6200 ;
      RECT 248.8500 0.0000 252.1500 0.6200 ;
      RECT 245.2500 0.0000 248.5500 0.6200 ;
      RECT 241.6500 0.0000 244.9500 0.6200 ;
      RECT 238.0500 0.0000 241.3500 0.6200 ;
      RECT 234.4500 0.0000 237.7500 0.6200 ;
      RECT 230.8500 0.0000 234.1500 0.6200 ;
      RECT 227.2500 0.0000 230.5500 0.6200 ;
      RECT 223.6500 0.0000 226.9500 0.6200 ;
      RECT 220.0500 0.0000 223.3500 0.6200 ;
      RECT 216.4500 0.0000 219.7500 0.6200 ;
      RECT 212.8500 0.0000 216.1500 0.6200 ;
      RECT 209.2500 0.0000 212.5500 0.6200 ;
      RECT 205.6500 0.0000 208.9500 0.6200 ;
      RECT 202.0500 0.0000 205.3500 0.6200 ;
      RECT 198.4500 0.0000 201.7500 0.6200 ;
      RECT 194.8500 0.0000 198.1500 0.6200 ;
      RECT 191.2500 0.0000 194.5500 0.6200 ;
      RECT 187.6500 0.0000 190.9500 0.6200 ;
      RECT 184.0500 0.0000 187.3500 0.6200 ;
      RECT 180.4500 0.0000 183.7500 0.6200 ;
      RECT 176.8500 0.0000 180.1500 0.6200 ;
      RECT 173.2500 0.0000 176.5500 0.6200 ;
      RECT 169.6500 0.0000 172.9500 0.6200 ;
      RECT 166.0500 0.0000 169.3500 0.6200 ;
      RECT 162.4500 0.0000 165.7500 0.6200 ;
      RECT 158.8500 0.0000 162.1500 0.6200 ;
      RECT 155.2500 0.0000 158.5500 0.6200 ;
      RECT 151.6500 0.0000 154.9500 0.6200 ;
      RECT 148.0500 0.0000 151.3500 0.6200 ;
      RECT 144.4500 0.0000 147.7500 0.6200 ;
      RECT 140.8500 0.0000 144.1500 0.6200 ;
      RECT 137.2500 0.0000 140.5500 0.6200 ;
      RECT 133.6500 0.0000 136.9500 0.6200 ;
      RECT 130.0500 0.0000 133.3500 0.6200 ;
      RECT 126.4500 0.0000 129.7500 0.6200 ;
      RECT 122.8500 0.0000 126.1500 0.6200 ;
      RECT 119.2500 0.0000 122.5500 0.6200 ;
      RECT 115.6500 0.0000 118.9500 0.6200 ;
      RECT 112.0500 0.0000 115.3500 0.6200 ;
      RECT 108.4500 0.0000 111.7500 0.6200 ;
      RECT 104.8500 0.0000 108.1500 0.6200 ;
      RECT 101.2500 0.0000 104.5500 0.6200 ;
      RECT 97.6500 0.0000 100.9500 0.6200 ;
      RECT 94.0500 0.0000 97.3500 0.6200 ;
      RECT 90.4500 0.0000 93.7500 0.6200 ;
      RECT 86.8500 0.0000 90.1500 0.6200 ;
      RECT 83.2500 0.0000 86.5500 0.6200 ;
      RECT 79.6500 0.0000 82.9500 0.6200 ;
      RECT 76.0500 0.0000 79.3500 0.6200 ;
      RECT 72.4500 0.0000 75.7500 0.6200 ;
      RECT 68.8500 0.0000 72.1500 0.6200 ;
      RECT 65.2500 0.0000 68.5500 0.6200 ;
      RECT 61.6500 0.0000 64.9500 0.6200 ;
      RECT 58.0500 0.0000 61.3500 0.6200 ;
      RECT 54.4500 0.0000 57.7500 0.6200 ;
      RECT 50.8500 0.0000 54.1500 0.6200 ;
      RECT 47.2500 0.0000 50.5500 0.6200 ;
      RECT 43.6500 0.0000 46.9500 0.6200 ;
      RECT 40.0500 0.0000 43.3500 0.6200 ;
      RECT 36.4500 0.0000 39.7500 0.6200 ;
      RECT 32.8500 0.0000 36.1500 0.6200 ;
      RECT 29.2500 0.0000 32.5500 0.6200 ;
      RECT 25.6500 0.0000 28.9500 0.6200 ;
      RECT 22.0500 0.0000 25.3500 0.6200 ;
      RECT 18.4500 0.0000 21.7500 0.6200 ;
      RECT 0.0000 0.0000 18.1500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 229.5500 608.8000 311.6000 ;
      RECT 0.6200 229.2500 608.8000 229.5500 ;
      RECT 0.0000 227.7500 608.8000 229.2500 ;
      RECT 0.6200 227.4500 608.8000 227.7500 ;
      RECT 0.0000 225.9500 608.8000 227.4500 ;
      RECT 0.6200 225.6500 608.8000 225.9500 ;
      RECT 0.0000 224.1500 608.8000 225.6500 ;
      RECT 0.6200 223.8500 608.8000 224.1500 ;
      RECT 0.0000 222.3500 608.8000 223.8500 ;
      RECT 0.6200 222.0500 608.8000 222.3500 ;
      RECT 0.0000 220.5500 608.8000 222.0500 ;
      RECT 0.6200 220.2500 608.8000 220.5500 ;
      RECT 0.0000 218.7500 608.8000 220.2500 ;
      RECT 0.6200 218.4500 608.8000 218.7500 ;
      RECT 0.0000 216.9500 608.8000 218.4500 ;
      RECT 0.6200 216.6500 608.8000 216.9500 ;
      RECT 0.0000 215.1500 608.8000 216.6500 ;
      RECT 0.6200 214.8500 608.8000 215.1500 ;
      RECT 0.0000 213.3500 608.8000 214.8500 ;
      RECT 0.6200 213.0500 608.8000 213.3500 ;
      RECT 0.0000 211.5500 608.8000 213.0500 ;
      RECT 0.6200 211.2500 608.8000 211.5500 ;
      RECT 0.0000 209.7500 608.8000 211.2500 ;
      RECT 0.6200 209.4500 608.8000 209.7500 ;
      RECT 0.0000 207.9500 608.8000 209.4500 ;
      RECT 0.6200 207.6500 608.8000 207.9500 ;
      RECT 0.0000 206.1500 608.8000 207.6500 ;
      RECT 0.6200 205.8500 608.8000 206.1500 ;
      RECT 0.0000 204.3500 608.8000 205.8500 ;
      RECT 0.6200 204.0500 608.8000 204.3500 ;
      RECT 0.0000 202.5500 608.8000 204.0500 ;
      RECT 0.6200 202.2500 608.8000 202.5500 ;
      RECT 0.0000 200.7500 608.8000 202.2500 ;
      RECT 0.6200 200.4500 608.8000 200.7500 ;
      RECT 0.0000 198.9500 608.8000 200.4500 ;
      RECT 0.6200 198.6500 608.8000 198.9500 ;
      RECT 0.0000 197.1500 608.8000 198.6500 ;
      RECT 0.6200 196.8500 608.8000 197.1500 ;
      RECT 0.0000 195.3500 608.8000 196.8500 ;
      RECT 0.6200 195.0500 608.8000 195.3500 ;
      RECT 0.0000 193.5500 608.8000 195.0500 ;
      RECT 0.6200 193.2500 608.8000 193.5500 ;
      RECT 0.0000 191.7500 608.8000 193.2500 ;
      RECT 0.6200 191.4500 608.8000 191.7500 ;
      RECT 0.0000 189.9500 608.8000 191.4500 ;
      RECT 0.6200 189.6500 608.8000 189.9500 ;
      RECT 0.0000 188.1500 608.8000 189.6500 ;
      RECT 0.6200 187.8500 608.8000 188.1500 ;
      RECT 0.0000 186.3500 608.8000 187.8500 ;
      RECT 0.6200 186.0500 608.8000 186.3500 ;
      RECT 0.0000 184.5500 608.8000 186.0500 ;
      RECT 0.6200 184.2500 608.8000 184.5500 ;
      RECT 0.0000 182.7500 608.8000 184.2500 ;
      RECT 0.6200 182.4500 608.8000 182.7500 ;
      RECT 0.0000 180.9500 608.8000 182.4500 ;
      RECT 0.6200 180.6500 608.8000 180.9500 ;
      RECT 0.0000 179.1500 608.8000 180.6500 ;
      RECT 0.6200 178.8500 608.8000 179.1500 ;
      RECT 0.0000 177.3500 608.8000 178.8500 ;
      RECT 0.6200 177.0500 608.8000 177.3500 ;
      RECT 0.0000 175.5500 608.8000 177.0500 ;
      RECT 0.6200 175.2500 608.8000 175.5500 ;
      RECT 0.0000 173.7500 608.8000 175.2500 ;
      RECT 0.6200 173.4500 608.8000 173.7500 ;
      RECT 0.0000 171.9500 608.8000 173.4500 ;
      RECT 0.6200 171.6500 608.8000 171.9500 ;
      RECT 0.0000 170.1500 608.8000 171.6500 ;
      RECT 0.6200 169.8500 608.8000 170.1500 ;
      RECT 0.0000 168.3500 608.8000 169.8500 ;
      RECT 0.6200 168.0500 608.8000 168.3500 ;
      RECT 0.0000 166.5500 608.8000 168.0500 ;
      RECT 0.6200 166.2500 608.8000 166.5500 ;
      RECT 0.0000 164.7500 608.8000 166.2500 ;
      RECT 0.6200 164.4500 608.8000 164.7500 ;
      RECT 0.0000 162.9500 608.8000 164.4500 ;
      RECT 0.6200 162.6500 608.8000 162.9500 ;
      RECT 0.0000 161.1500 608.8000 162.6500 ;
      RECT 0.6200 160.8500 608.8000 161.1500 ;
      RECT 0.0000 159.3500 608.8000 160.8500 ;
      RECT 0.6200 159.0500 608.8000 159.3500 ;
      RECT 0.0000 157.5500 608.8000 159.0500 ;
      RECT 0.6200 157.2500 608.8000 157.5500 ;
      RECT 0.0000 155.7500 608.8000 157.2500 ;
      RECT 0.6200 155.4500 608.8000 155.7500 ;
      RECT 0.0000 153.9500 608.8000 155.4500 ;
      RECT 0.6200 153.6500 608.8000 153.9500 ;
      RECT 0.0000 152.1500 608.8000 153.6500 ;
      RECT 0.6200 151.8500 608.8000 152.1500 ;
      RECT 0.0000 150.3500 608.8000 151.8500 ;
      RECT 0.6200 150.0500 608.8000 150.3500 ;
      RECT 0.0000 148.5500 608.8000 150.0500 ;
      RECT 0.6200 148.2500 608.8000 148.5500 ;
      RECT 0.0000 146.7500 608.8000 148.2500 ;
      RECT 0.6200 146.4500 608.8000 146.7500 ;
      RECT 0.0000 144.9500 608.8000 146.4500 ;
      RECT 0.6200 144.6500 608.8000 144.9500 ;
      RECT 0.0000 143.1500 608.8000 144.6500 ;
      RECT 0.6200 142.8500 608.8000 143.1500 ;
      RECT 0.0000 141.3500 608.8000 142.8500 ;
      RECT 0.6200 141.0500 608.8000 141.3500 ;
      RECT 0.0000 139.5500 608.8000 141.0500 ;
      RECT 0.6200 139.2500 608.8000 139.5500 ;
      RECT 0.0000 137.7500 608.8000 139.2500 ;
      RECT 0.6200 137.4500 608.8000 137.7500 ;
      RECT 0.0000 135.9500 608.8000 137.4500 ;
      RECT 0.6200 135.6500 608.8000 135.9500 ;
      RECT 0.0000 134.1500 608.8000 135.6500 ;
      RECT 0.6200 133.8500 608.8000 134.1500 ;
      RECT 0.0000 132.3500 608.8000 133.8500 ;
      RECT 0.6200 132.0500 608.8000 132.3500 ;
      RECT 0.0000 130.5500 608.8000 132.0500 ;
      RECT 0.6200 130.2500 608.8000 130.5500 ;
      RECT 0.0000 128.7500 608.8000 130.2500 ;
      RECT 0.6200 128.4500 608.8000 128.7500 ;
      RECT 0.0000 126.9500 608.8000 128.4500 ;
      RECT 0.6200 126.6500 608.8000 126.9500 ;
      RECT 0.0000 125.1500 608.8000 126.6500 ;
      RECT 0.6200 124.8500 608.8000 125.1500 ;
      RECT 0.0000 123.3500 608.8000 124.8500 ;
      RECT 0.6200 123.0500 608.8000 123.3500 ;
      RECT 0.0000 121.5500 608.8000 123.0500 ;
      RECT 0.6200 121.2500 608.8000 121.5500 ;
      RECT 0.0000 119.7500 608.8000 121.2500 ;
      RECT 0.6200 119.4500 608.8000 119.7500 ;
      RECT 0.0000 117.9500 608.8000 119.4500 ;
      RECT 0.6200 117.6500 608.8000 117.9500 ;
      RECT 0.0000 116.1500 608.8000 117.6500 ;
      RECT 0.6200 115.8500 608.8000 116.1500 ;
      RECT 0.0000 114.3500 608.8000 115.8500 ;
      RECT 0.6200 114.0500 608.8000 114.3500 ;
      RECT 0.0000 112.5500 608.8000 114.0500 ;
      RECT 0.6200 112.2500 608.8000 112.5500 ;
      RECT 0.0000 110.7500 608.8000 112.2500 ;
      RECT 0.6200 110.4500 608.8000 110.7500 ;
      RECT 0.0000 108.9500 608.8000 110.4500 ;
      RECT 0.6200 108.6500 608.8000 108.9500 ;
      RECT 0.0000 107.1500 608.8000 108.6500 ;
      RECT 0.6200 106.8500 608.8000 107.1500 ;
      RECT 0.0000 105.3500 608.8000 106.8500 ;
      RECT 0.6200 105.0500 608.8000 105.3500 ;
      RECT 0.0000 103.5500 608.8000 105.0500 ;
      RECT 0.6200 103.2500 608.8000 103.5500 ;
      RECT 0.0000 101.7500 608.8000 103.2500 ;
      RECT 0.6200 101.4500 608.8000 101.7500 ;
      RECT 0.0000 99.9500 608.8000 101.4500 ;
      RECT 0.6200 99.6500 608.8000 99.9500 ;
      RECT 0.0000 98.1500 608.8000 99.6500 ;
      RECT 0.6200 97.8500 608.8000 98.1500 ;
      RECT 0.0000 96.3500 608.8000 97.8500 ;
      RECT 0.6200 96.0500 608.8000 96.3500 ;
      RECT 0.0000 94.5500 608.8000 96.0500 ;
      RECT 0.6200 94.2500 608.8000 94.5500 ;
      RECT 0.0000 92.7500 608.8000 94.2500 ;
      RECT 0.6200 92.4500 608.8000 92.7500 ;
      RECT 0.0000 90.9500 608.8000 92.4500 ;
      RECT 0.6200 90.6500 608.8000 90.9500 ;
      RECT 0.0000 89.1500 608.8000 90.6500 ;
      RECT 0.6200 88.8500 608.8000 89.1500 ;
      RECT 0.0000 87.3500 608.8000 88.8500 ;
      RECT 0.6200 87.0500 608.8000 87.3500 ;
      RECT 0.0000 85.5500 608.8000 87.0500 ;
      RECT 0.6200 85.2500 608.8000 85.5500 ;
      RECT 0.0000 83.7500 608.8000 85.2500 ;
      RECT 0.6200 83.4500 608.8000 83.7500 ;
      RECT 0.0000 81.9500 608.8000 83.4500 ;
      RECT 0.6200 81.6500 608.8000 81.9500 ;
      RECT 0.0000 0.0000 608.8000 81.6500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 608.8000 311.6000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 608.8000 311.6000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 608.8000 311.6000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 608.8000 311.6000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 608.8000 311.6000 ;
  END
END core

END LIBRARY
