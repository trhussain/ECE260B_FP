/home/linux/ieng6/ee260bwi25/aekeng/ECE260B_FP/ece260_project/step3/pnr/pnrTopModule/subckt/sram_w16_160.lef