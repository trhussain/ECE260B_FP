/home/linux/ieng6/ee260bwi25/aekeng/test/ECE260B_FP/ece260_project/step3/pnr2/subckt/sram_w16_64.lef