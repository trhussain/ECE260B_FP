##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 22 17:45:17 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 381.2000 BY 380.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 1.1500 0.5200 1.2500 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 243.3500 0.5200 243.4500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 240.3500 0.5200 240.4500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 237.3500 0.5200 237.4500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 234.3500 0.5200 234.4500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 231.3500 0.5200 231.4500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 228.3500 0.5200 228.4500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 225.3500 0.5200 225.4500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 222.3500 0.5200 222.4500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 219.3500 0.5200 219.4500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 216.3500 0.5200 216.4500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 213.3500 0.5200 213.4500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 210.3500 0.5200 210.4500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 207.3500 0.5200 207.4500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 204.3500 0.5200 204.4500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 201.3500 0.5200 201.4500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 198.3500 0.5200 198.4500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 195.3500 0.5200 195.4500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 192.3500 0.5200 192.4500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 189.3500 0.5200 189.4500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 186.3500 0.5200 186.4500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 183.3500 0.5200 183.4500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 180.3500 0.5200 180.4500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 177.3500 0.5200 177.4500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 174.3500 0.5200 174.4500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 171.3500 0.5200 171.4500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 168.3500 0.5200 168.4500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 165.3500 0.5200 165.4500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 162.3500 0.5200 162.4500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 159.3500 0.5200 159.4500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 156.3500 0.5200 156.4500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 153.3500 0.5200 153.4500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 150.3500 0.5200 150.4500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 147.3500 0.5200 147.4500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 144.3500 0.5200 144.4500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 141.3500 0.5200 141.4500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 138.3500 0.5200 138.4500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 135.3500 0.5200 135.4500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 132.3500 0.5200 132.4500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 129.3500 0.5200 129.4500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 126.3500 0.5200 126.4500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 123.3500 0.5200 123.4500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 120.3500 0.5200 120.4500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 117.3500 0.5200 117.4500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 114.3500 0.5200 114.4500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 111.3500 0.5200 111.4500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 108.3500 0.5200 108.4500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 105.3500 0.5200 105.4500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 102.3500 0.5200 102.4500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 99.3500 0.5200 99.4500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 96.3500 0.5200 96.4500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 93.3500 0.5200 93.4500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 90.3500 0.5200 90.4500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 87.3500 0.5200 87.4500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 84.3500 0.5200 84.4500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 81.3500 0.5200 81.4500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 78.3500 0.5200 78.4500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 75.3500 0.5200 75.4500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 72.3500 0.5200 72.4500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 69.3500 0.5200 69.4500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 66.3500 0.5200 66.4500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 63.3500 0.5200 63.4500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 60.3500 0.5200 60.4500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.3500 0.5200 57.4500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 54.3500 0.5200 54.4500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.2500 0.0000 34.3500 0.5200 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.2500 0.0000 36.3500 0.5200 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.2500 0.0000 38.3500 0.5200 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.2500 0.0000 40.3500 0.5200 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.2500 0.0000 42.3500 0.5200 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.2500 0.0000 44.3500 0.5200 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.2500 0.0000 46.3500 0.5200 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.2500 0.0000 48.3500 0.5200 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.2500 0.0000 50.3500 0.5200 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.2500 0.0000 52.3500 0.5200 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.2500 0.0000 54.3500 0.5200 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.2500 0.0000 56.3500 0.5200 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.2500 0.0000 58.3500 0.5200 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.2500 0.0000 60.3500 0.5200 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.2500 0.0000 62.3500 0.5200 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.2500 0.0000 64.3500 0.5200 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.2500 0.0000 66.3500 0.5200 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.2500 0.0000 68.3500 0.5200 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.2500 0.0000 70.3500 0.5200 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.2500 0.0000 72.3500 0.5200 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.2500 0.0000 74.3500 0.5200 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.2500 0.0000 76.3500 0.5200 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.2500 0.0000 78.3500 0.5200 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.2500 0.0000 80.3500 0.5200 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.2500 0.0000 82.3500 0.5200 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.2500 0.0000 84.3500 0.5200 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.2500 0.0000 86.3500 0.5200 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.2500 0.0000 88.3500 0.5200 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.2500 0.0000 90.3500 0.5200 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.2500 0.0000 92.3500 0.5200 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.2500 0.0000 94.3500 0.5200 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.2500 0.0000 96.3500 0.5200 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.2500 0.0000 98.3500 0.5200 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.2500 0.0000 100.3500 0.5200 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.2500 0.0000 102.3500 0.5200 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.2500 0.0000 104.3500 0.5200 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.2500 0.0000 106.3500 0.5200 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.2500 0.0000 108.3500 0.5200 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.2500 0.0000 110.3500 0.5200 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.2500 0.0000 112.3500 0.5200 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.2500 0.0000 114.3500 0.5200 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.2500 0.0000 116.3500 0.5200 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.2500 0.0000 118.3500 0.5200 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.2500 0.0000 120.3500 0.5200 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.2500 0.0000 122.3500 0.5200 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.2500 0.0000 124.3500 0.5200 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.2500 0.0000 126.3500 0.5200 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.2500 0.0000 128.3500 0.5200 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.2500 0.0000 130.3500 0.5200 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.2500 0.0000 132.3500 0.5200 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.2500 0.0000 134.3500 0.5200 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.2500 0.0000 136.3500 0.5200 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.2500 0.0000 138.3500 0.5200 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.2500 0.0000 140.3500 0.5200 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.2500 0.0000 142.3500 0.5200 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.2500 0.0000 144.3500 0.5200 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.2500 0.0000 146.3500 0.5200 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.2500 0.0000 148.3500 0.5200 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.2500 0.0000 150.3500 0.5200 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.2500 0.0000 152.3500 0.5200 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.2500 0.0000 154.3500 0.5200 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.2500 0.0000 156.3500 0.5200 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.2500 0.0000 158.3500 0.5200 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.2500 0.0000 160.3500 0.5200 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.2500 0.0000 162.3500 0.5200 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.2500 0.0000 164.3500 0.5200 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.2500 0.0000 166.3500 0.5200 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.2500 0.0000 168.3500 0.5200 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.2500 0.0000 170.3500 0.5200 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.2500 0.0000 172.3500 0.5200 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.2500 0.0000 174.3500 0.5200 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.2500 0.0000 176.3500 0.5200 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.2500 0.0000 178.3500 0.5200 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.2500 0.0000 180.3500 0.5200 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.2500 0.0000 182.3500 0.5200 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.2500 0.0000 184.3500 0.5200 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.2500 0.0000 186.3500 0.5200 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.2500 0.0000 188.3500 0.5200 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.2500 0.0000 190.3500 0.5200 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.2500 0.0000 192.3500 0.5200 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.2500 0.0000 194.3500 0.5200 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.2500 0.0000 196.3500 0.5200 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.2500 0.0000 198.3500 0.5200 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.2500 0.0000 200.3500 0.5200 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.2500 0.0000 202.3500 0.5200 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.2500 0.0000 204.3500 0.5200 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 206.2500 0.0000 206.3500 0.5200 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.2500 0.0000 208.3500 0.5200 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.2500 0.0000 210.3500 0.5200 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.2500 0.0000 212.3500 0.5200 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.2500 0.0000 214.3500 0.5200 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.2500 0.0000 216.3500 0.5200 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.2500 0.0000 218.3500 0.5200 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.2500 0.0000 220.3500 0.5200 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.2500 0.0000 222.3500 0.5200 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.2500 0.0000 224.3500 0.5200 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.2500 0.0000 226.3500 0.5200 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.2500 0.0000 228.3500 0.5200 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.2500 0.0000 230.3500 0.5200 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.2500 0.0000 232.3500 0.5200 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.2500 0.0000 234.3500 0.5200 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 236.2500 0.0000 236.3500 0.5200 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.2500 0.0000 238.3500 0.5200 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.2500 0.0000 240.3500 0.5200 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 242.2500 0.0000 242.3500 0.5200 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 244.2500 0.0000 244.3500 0.5200 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.2500 0.0000 246.3500 0.5200 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.2500 0.0000 248.3500 0.5200 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 250.2500 0.0000 250.3500 0.5200 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.2500 0.0000 252.3500 0.5200 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 254.2500 0.0000 254.3500 0.5200 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.2500 0.0000 256.3500 0.5200 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 258.2500 0.0000 258.3500 0.5200 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.2500 0.0000 260.3500 0.5200 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.2500 0.0000 262.3500 0.5200 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 264.2500 0.0000 264.3500 0.5200 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 266.2500 0.0000 266.3500 0.5200 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 268.2500 0.0000 268.3500 0.5200 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.2500 0.0000 270.3500 0.5200 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 272.2500 0.0000 272.3500 0.5200 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.2500 0.0000 274.3500 0.5200 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 276.2500 0.0000 276.3500 0.5200 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.2500 0.0000 278.3500 0.5200 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.2500 0.0000 280.3500 0.5200 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.2500 0.0000 282.3500 0.5200 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284.2500 0.0000 284.3500 0.5200 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 286.2500 0.0000 286.3500 0.5200 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.2500 0.0000 288.3500 0.5200 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 290.2500 0.0000 290.3500 0.5200 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 292.2500 0.0000 292.3500 0.5200 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 294.2500 0.0000 294.3500 0.5200 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 296.2500 0.0000 296.3500 0.5200 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 298.2500 0.0000 298.3500 0.5200 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.2500 0.0000 300.3500 0.5200 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.2500 0.0000 302.3500 0.5200 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 304.2500 0.0000 304.3500 0.5200 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.2500 0.0000 306.3500 0.5200 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.2500 0.0000 308.3500 0.5200 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.2500 0.0000 310.3500 0.5200 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.2500 0.0000 312.3500 0.5200 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.2500 0.0000 314.3500 0.5200 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.2500 0.0000 316.3500 0.5200 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.2500 0.0000 318.3500 0.5200 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.2500 0.0000 320.3500 0.5200 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.2500 0.0000 322.3500 0.5200 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.2500 0.0000 324.3500 0.5200 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.2500 0.0000 326.3500 0.5200 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.2500 0.0000 328.3500 0.5200 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.2500 0.0000 330.3500 0.5200 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.2500 0.0000 332.3500 0.5200 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.2500 0.0000 334.3500 0.5200 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.2500 0.0000 336.3500 0.5200 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.2500 0.0000 338.3500 0.5200 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.2500 0.0000 340.3500 0.5200 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.2500 0.0000 342.3500 0.5200 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.2500 0.0000 344.3500 0.5200 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.2500 0.0000 346.3500 0.5200 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.2500 0.0000 348.3500 0.5200 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.2500 0.0000 350.3500 0.5200 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.2500 0.0000 352.3500 0.5200 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 51.3500 0.5200 51.4500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 48.3500 0.5200 48.4500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 45.3500 0.5200 45.4500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 42.3500 0.5200 42.4500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 39.3500 0.5200 39.4500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.3500 0.5200 36.4500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.3500 0.5200 33.4500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.3500 0.5200 30.4500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.3500 0.5200 27.4500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.3500 0.5200 24.4500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.3500 0.5200 21.4500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.3500 0.5200 18.4500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.3500 0.5200 15.4500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 12.3500 0.5200 12.4500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 9.3500 0.5200 9.4500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 6.3500 0.5200 6.4500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 3.3500 0.5200 3.4500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 246.3500 0.5200 246.4500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 381.2000 380.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.6200 381.2000 380.0000 ;
      RECT 352.4500 0.0000 381.2000 0.6200 ;
      RECT 350.4500 0.0000 352.1500 0.6200 ;
      RECT 348.4500 0.0000 350.1500 0.6200 ;
      RECT 346.4500 0.0000 348.1500 0.6200 ;
      RECT 344.4500 0.0000 346.1500 0.6200 ;
      RECT 342.4500 0.0000 344.1500 0.6200 ;
      RECT 340.4500 0.0000 342.1500 0.6200 ;
      RECT 338.4500 0.0000 340.1500 0.6200 ;
      RECT 336.4500 0.0000 338.1500 0.6200 ;
      RECT 334.4500 0.0000 336.1500 0.6200 ;
      RECT 332.4500 0.0000 334.1500 0.6200 ;
      RECT 330.4500 0.0000 332.1500 0.6200 ;
      RECT 328.4500 0.0000 330.1500 0.6200 ;
      RECT 326.4500 0.0000 328.1500 0.6200 ;
      RECT 324.4500 0.0000 326.1500 0.6200 ;
      RECT 322.4500 0.0000 324.1500 0.6200 ;
      RECT 320.4500 0.0000 322.1500 0.6200 ;
      RECT 318.4500 0.0000 320.1500 0.6200 ;
      RECT 316.4500 0.0000 318.1500 0.6200 ;
      RECT 314.4500 0.0000 316.1500 0.6200 ;
      RECT 312.4500 0.0000 314.1500 0.6200 ;
      RECT 310.4500 0.0000 312.1500 0.6200 ;
      RECT 308.4500 0.0000 310.1500 0.6200 ;
      RECT 306.4500 0.0000 308.1500 0.6200 ;
      RECT 304.4500 0.0000 306.1500 0.6200 ;
      RECT 302.4500 0.0000 304.1500 0.6200 ;
      RECT 300.4500 0.0000 302.1500 0.6200 ;
      RECT 298.4500 0.0000 300.1500 0.6200 ;
      RECT 296.4500 0.0000 298.1500 0.6200 ;
      RECT 294.4500 0.0000 296.1500 0.6200 ;
      RECT 292.4500 0.0000 294.1500 0.6200 ;
      RECT 290.4500 0.0000 292.1500 0.6200 ;
      RECT 288.4500 0.0000 290.1500 0.6200 ;
      RECT 286.4500 0.0000 288.1500 0.6200 ;
      RECT 284.4500 0.0000 286.1500 0.6200 ;
      RECT 282.4500 0.0000 284.1500 0.6200 ;
      RECT 280.4500 0.0000 282.1500 0.6200 ;
      RECT 278.4500 0.0000 280.1500 0.6200 ;
      RECT 276.4500 0.0000 278.1500 0.6200 ;
      RECT 274.4500 0.0000 276.1500 0.6200 ;
      RECT 272.4500 0.0000 274.1500 0.6200 ;
      RECT 270.4500 0.0000 272.1500 0.6200 ;
      RECT 268.4500 0.0000 270.1500 0.6200 ;
      RECT 266.4500 0.0000 268.1500 0.6200 ;
      RECT 264.4500 0.0000 266.1500 0.6200 ;
      RECT 262.4500 0.0000 264.1500 0.6200 ;
      RECT 260.4500 0.0000 262.1500 0.6200 ;
      RECT 258.4500 0.0000 260.1500 0.6200 ;
      RECT 256.4500 0.0000 258.1500 0.6200 ;
      RECT 254.4500 0.0000 256.1500 0.6200 ;
      RECT 252.4500 0.0000 254.1500 0.6200 ;
      RECT 250.4500 0.0000 252.1500 0.6200 ;
      RECT 248.4500 0.0000 250.1500 0.6200 ;
      RECT 246.4500 0.0000 248.1500 0.6200 ;
      RECT 244.4500 0.0000 246.1500 0.6200 ;
      RECT 242.4500 0.0000 244.1500 0.6200 ;
      RECT 240.4500 0.0000 242.1500 0.6200 ;
      RECT 238.4500 0.0000 240.1500 0.6200 ;
      RECT 236.4500 0.0000 238.1500 0.6200 ;
      RECT 234.4500 0.0000 236.1500 0.6200 ;
      RECT 232.4500 0.0000 234.1500 0.6200 ;
      RECT 230.4500 0.0000 232.1500 0.6200 ;
      RECT 228.4500 0.0000 230.1500 0.6200 ;
      RECT 226.4500 0.0000 228.1500 0.6200 ;
      RECT 224.4500 0.0000 226.1500 0.6200 ;
      RECT 222.4500 0.0000 224.1500 0.6200 ;
      RECT 220.4500 0.0000 222.1500 0.6200 ;
      RECT 218.4500 0.0000 220.1500 0.6200 ;
      RECT 216.4500 0.0000 218.1500 0.6200 ;
      RECT 214.4500 0.0000 216.1500 0.6200 ;
      RECT 212.4500 0.0000 214.1500 0.6200 ;
      RECT 210.4500 0.0000 212.1500 0.6200 ;
      RECT 208.4500 0.0000 210.1500 0.6200 ;
      RECT 206.4500 0.0000 208.1500 0.6200 ;
      RECT 204.4500 0.0000 206.1500 0.6200 ;
      RECT 202.4500 0.0000 204.1500 0.6200 ;
      RECT 200.4500 0.0000 202.1500 0.6200 ;
      RECT 198.4500 0.0000 200.1500 0.6200 ;
      RECT 196.4500 0.0000 198.1500 0.6200 ;
      RECT 194.4500 0.0000 196.1500 0.6200 ;
      RECT 192.4500 0.0000 194.1500 0.6200 ;
      RECT 190.4500 0.0000 192.1500 0.6200 ;
      RECT 188.4500 0.0000 190.1500 0.6200 ;
      RECT 186.4500 0.0000 188.1500 0.6200 ;
      RECT 184.4500 0.0000 186.1500 0.6200 ;
      RECT 182.4500 0.0000 184.1500 0.6200 ;
      RECT 180.4500 0.0000 182.1500 0.6200 ;
      RECT 178.4500 0.0000 180.1500 0.6200 ;
      RECT 176.4500 0.0000 178.1500 0.6200 ;
      RECT 174.4500 0.0000 176.1500 0.6200 ;
      RECT 172.4500 0.0000 174.1500 0.6200 ;
      RECT 170.4500 0.0000 172.1500 0.6200 ;
      RECT 168.4500 0.0000 170.1500 0.6200 ;
      RECT 166.4500 0.0000 168.1500 0.6200 ;
      RECT 164.4500 0.0000 166.1500 0.6200 ;
      RECT 162.4500 0.0000 164.1500 0.6200 ;
      RECT 160.4500 0.0000 162.1500 0.6200 ;
      RECT 158.4500 0.0000 160.1500 0.6200 ;
      RECT 156.4500 0.0000 158.1500 0.6200 ;
      RECT 154.4500 0.0000 156.1500 0.6200 ;
      RECT 152.4500 0.0000 154.1500 0.6200 ;
      RECT 150.4500 0.0000 152.1500 0.6200 ;
      RECT 148.4500 0.0000 150.1500 0.6200 ;
      RECT 146.4500 0.0000 148.1500 0.6200 ;
      RECT 144.4500 0.0000 146.1500 0.6200 ;
      RECT 142.4500 0.0000 144.1500 0.6200 ;
      RECT 140.4500 0.0000 142.1500 0.6200 ;
      RECT 138.4500 0.0000 140.1500 0.6200 ;
      RECT 136.4500 0.0000 138.1500 0.6200 ;
      RECT 134.4500 0.0000 136.1500 0.6200 ;
      RECT 132.4500 0.0000 134.1500 0.6200 ;
      RECT 130.4500 0.0000 132.1500 0.6200 ;
      RECT 128.4500 0.0000 130.1500 0.6200 ;
      RECT 126.4500 0.0000 128.1500 0.6200 ;
      RECT 124.4500 0.0000 126.1500 0.6200 ;
      RECT 122.4500 0.0000 124.1500 0.6200 ;
      RECT 120.4500 0.0000 122.1500 0.6200 ;
      RECT 118.4500 0.0000 120.1500 0.6200 ;
      RECT 116.4500 0.0000 118.1500 0.6200 ;
      RECT 114.4500 0.0000 116.1500 0.6200 ;
      RECT 112.4500 0.0000 114.1500 0.6200 ;
      RECT 110.4500 0.0000 112.1500 0.6200 ;
      RECT 108.4500 0.0000 110.1500 0.6200 ;
      RECT 106.4500 0.0000 108.1500 0.6200 ;
      RECT 104.4500 0.0000 106.1500 0.6200 ;
      RECT 102.4500 0.0000 104.1500 0.6200 ;
      RECT 100.4500 0.0000 102.1500 0.6200 ;
      RECT 98.4500 0.0000 100.1500 0.6200 ;
      RECT 96.4500 0.0000 98.1500 0.6200 ;
      RECT 94.4500 0.0000 96.1500 0.6200 ;
      RECT 92.4500 0.0000 94.1500 0.6200 ;
      RECT 90.4500 0.0000 92.1500 0.6200 ;
      RECT 88.4500 0.0000 90.1500 0.6200 ;
      RECT 86.4500 0.0000 88.1500 0.6200 ;
      RECT 84.4500 0.0000 86.1500 0.6200 ;
      RECT 82.4500 0.0000 84.1500 0.6200 ;
      RECT 80.4500 0.0000 82.1500 0.6200 ;
      RECT 78.4500 0.0000 80.1500 0.6200 ;
      RECT 76.4500 0.0000 78.1500 0.6200 ;
      RECT 74.4500 0.0000 76.1500 0.6200 ;
      RECT 72.4500 0.0000 74.1500 0.6200 ;
      RECT 70.4500 0.0000 72.1500 0.6200 ;
      RECT 68.4500 0.0000 70.1500 0.6200 ;
      RECT 66.4500 0.0000 68.1500 0.6200 ;
      RECT 64.4500 0.0000 66.1500 0.6200 ;
      RECT 62.4500 0.0000 64.1500 0.6200 ;
      RECT 60.4500 0.0000 62.1500 0.6200 ;
      RECT 58.4500 0.0000 60.1500 0.6200 ;
      RECT 56.4500 0.0000 58.1500 0.6200 ;
      RECT 54.4500 0.0000 56.1500 0.6200 ;
      RECT 52.4500 0.0000 54.1500 0.6200 ;
      RECT 50.4500 0.0000 52.1500 0.6200 ;
      RECT 48.4500 0.0000 50.1500 0.6200 ;
      RECT 46.4500 0.0000 48.1500 0.6200 ;
      RECT 44.4500 0.0000 46.1500 0.6200 ;
      RECT 42.4500 0.0000 44.1500 0.6200 ;
      RECT 40.4500 0.0000 42.1500 0.6200 ;
      RECT 38.4500 0.0000 40.1500 0.6200 ;
      RECT 36.4500 0.0000 38.1500 0.6200 ;
      RECT 34.4500 0.0000 36.1500 0.6200 ;
      RECT 0.0000 0.0000 34.1500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 246.5500 381.2000 380.0000 ;
      RECT 0.6200 246.2500 381.2000 246.5500 ;
      RECT 0.0000 243.5500 381.2000 246.2500 ;
      RECT 0.6200 243.2500 381.2000 243.5500 ;
      RECT 0.0000 240.5500 381.2000 243.2500 ;
      RECT 0.6200 240.2500 381.2000 240.5500 ;
      RECT 0.0000 237.5500 381.2000 240.2500 ;
      RECT 0.6200 237.2500 381.2000 237.5500 ;
      RECT 0.0000 234.5500 381.2000 237.2500 ;
      RECT 0.6200 234.2500 381.2000 234.5500 ;
      RECT 0.0000 231.5500 381.2000 234.2500 ;
      RECT 0.6200 231.2500 381.2000 231.5500 ;
      RECT 0.0000 228.5500 381.2000 231.2500 ;
      RECT 0.6200 228.2500 381.2000 228.5500 ;
      RECT 0.0000 225.5500 381.2000 228.2500 ;
      RECT 0.6200 225.2500 381.2000 225.5500 ;
      RECT 0.0000 222.5500 381.2000 225.2500 ;
      RECT 0.6200 222.2500 381.2000 222.5500 ;
      RECT 0.0000 219.5500 381.2000 222.2500 ;
      RECT 0.6200 219.2500 381.2000 219.5500 ;
      RECT 0.0000 216.5500 381.2000 219.2500 ;
      RECT 0.6200 216.2500 381.2000 216.5500 ;
      RECT 0.0000 213.5500 381.2000 216.2500 ;
      RECT 0.6200 213.2500 381.2000 213.5500 ;
      RECT 0.0000 210.5500 381.2000 213.2500 ;
      RECT 0.6200 210.2500 381.2000 210.5500 ;
      RECT 0.0000 207.5500 381.2000 210.2500 ;
      RECT 0.6200 207.2500 381.2000 207.5500 ;
      RECT 0.0000 204.5500 381.2000 207.2500 ;
      RECT 0.6200 204.2500 381.2000 204.5500 ;
      RECT 0.0000 201.5500 381.2000 204.2500 ;
      RECT 0.6200 201.2500 381.2000 201.5500 ;
      RECT 0.0000 198.5500 381.2000 201.2500 ;
      RECT 0.6200 198.2500 381.2000 198.5500 ;
      RECT 0.0000 195.5500 381.2000 198.2500 ;
      RECT 0.6200 195.2500 381.2000 195.5500 ;
      RECT 0.0000 192.5500 381.2000 195.2500 ;
      RECT 0.6200 192.2500 381.2000 192.5500 ;
      RECT 0.0000 189.5500 381.2000 192.2500 ;
      RECT 0.6200 189.2500 381.2000 189.5500 ;
      RECT 0.0000 186.5500 381.2000 189.2500 ;
      RECT 0.6200 186.2500 381.2000 186.5500 ;
      RECT 0.0000 183.5500 381.2000 186.2500 ;
      RECT 0.6200 183.2500 381.2000 183.5500 ;
      RECT 0.0000 180.5500 381.2000 183.2500 ;
      RECT 0.6200 180.2500 381.2000 180.5500 ;
      RECT 0.0000 177.5500 381.2000 180.2500 ;
      RECT 0.6200 177.2500 381.2000 177.5500 ;
      RECT 0.0000 174.5500 381.2000 177.2500 ;
      RECT 0.6200 174.2500 381.2000 174.5500 ;
      RECT 0.0000 171.5500 381.2000 174.2500 ;
      RECT 0.6200 171.2500 381.2000 171.5500 ;
      RECT 0.0000 168.5500 381.2000 171.2500 ;
      RECT 0.6200 168.2500 381.2000 168.5500 ;
      RECT 0.0000 165.5500 381.2000 168.2500 ;
      RECT 0.6200 165.2500 381.2000 165.5500 ;
      RECT 0.0000 162.5500 381.2000 165.2500 ;
      RECT 0.6200 162.2500 381.2000 162.5500 ;
      RECT 0.0000 159.5500 381.2000 162.2500 ;
      RECT 0.6200 159.2500 381.2000 159.5500 ;
      RECT 0.0000 156.5500 381.2000 159.2500 ;
      RECT 0.6200 156.2500 381.2000 156.5500 ;
      RECT 0.0000 153.5500 381.2000 156.2500 ;
      RECT 0.6200 153.2500 381.2000 153.5500 ;
      RECT 0.0000 150.5500 381.2000 153.2500 ;
      RECT 0.6200 150.2500 381.2000 150.5500 ;
      RECT 0.0000 147.5500 381.2000 150.2500 ;
      RECT 0.6200 147.2500 381.2000 147.5500 ;
      RECT 0.0000 144.5500 381.2000 147.2500 ;
      RECT 0.6200 144.2500 381.2000 144.5500 ;
      RECT 0.0000 141.5500 381.2000 144.2500 ;
      RECT 0.6200 141.2500 381.2000 141.5500 ;
      RECT 0.0000 138.5500 381.2000 141.2500 ;
      RECT 0.6200 138.2500 381.2000 138.5500 ;
      RECT 0.0000 135.5500 381.2000 138.2500 ;
      RECT 0.6200 135.2500 381.2000 135.5500 ;
      RECT 0.0000 132.5500 381.2000 135.2500 ;
      RECT 0.6200 132.2500 381.2000 132.5500 ;
      RECT 0.0000 129.5500 381.2000 132.2500 ;
      RECT 0.6200 129.2500 381.2000 129.5500 ;
      RECT 0.0000 126.5500 381.2000 129.2500 ;
      RECT 0.6200 126.2500 381.2000 126.5500 ;
      RECT 0.0000 123.5500 381.2000 126.2500 ;
      RECT 0.6200 123.2500 381.2000 123.5500 ;
      RECT 0.0000 120.5500 381.2000 123.2500 ;
      RECT 0.6200 120.2500 381.2000 120.5500 ;
      RECT 0.0000 117.5500 381.2000 120.2500 ;
      RECT 0.6200 117.2500 381.2000 117.5500 ;
      RECT 0.0000 114.5500 381.2000 117.2500 ;
      RECT 0.6200 114.2500 381.2000 114.5500 ;
      RECT 0.0000 111.5500 381.2000 114.2500 ;
      RECT 0.6200 111.2500 381.2000 111.5500 ;
      RECT 0.0000 108.5500 381.2000 111.2500 ;
      RECT 0.6200 108.2500 381.2000 108.5500 ;
      RECT 0.0000 105.5500 381.2000 108.2500 ;
      RECT 0.6200 105.2500 381.2000 105.5500 ;
      RECT 0.0000 102.5500 381.2000 105.2500 ;
      RECT 0.6200 102.2500 381.2000 102.5500 ;
      RECT 0.0000 99.5500 381.2000 102.2500 ;
      RECT 0.6200 99.2500 381.2000 99.5500 ;
      RECT 0.0000 96.5500 381.2000 99.2500 ;
      RECT 0.6200 96.2500 381.2000 96.5500 ;
      RECT 0.0000 93.5500 381.2000 96.2500 ;
      RECT 0.6200 93.2500 381.2000 93.5500 ;
      RECT 0.0000 90.5500 381.2000 93.2500 ;
      RECT 0.6200 90.2500 381.2000 90.5500 ;
      RECT 0.0000 87.5500 381.2000 90.2500 ;
      RECT 0.6200 87.2500 381.2000 87.5500 ;
      RECT 0.0000 84.5500 381.2000 87.2500 ;
      RECT 0.6200 84.2500 381.2000 84.5500 ;
      RECT 0.0000 81.5500 381.2000 84.2500 ;
      RECT 0.6200 81.2500 381.2000 81.5500 ;
      RECT 0.0000 78.5500 381.2000 81.2500 ;
      RECT 0.6200 78.2500 381.2000 78.5500 ;
      RECT 0.0000 75.5500 381.2000 78.2500 ;
      RECT 0.6200 75.2500 381.2000 75.5500 ;
      RECT 0.0000 72.5500 381.2000 75.2500 ;
      RECT 0.6200 72.2500 381.2000 72.5500 ;
      RECT 0.0000 69.5500 381.2000 72.2500 ;
      RECT 0.6200 69.2500 381.2000 69.5500 ;
      RECT 0.0000 66.5500 381.2000 69.2500 ;
      RECT 0.6200 66.2500 381.2000 66.5500 ;
      RECT 0.0000 63.5500 381.2000 66.2500 ;
      RECT 0.6200 63.2500 381.2000 63.5500 ;
      RECT 0.0000 60.5500 381.2000 63.2500 ;
      RECT 0.6200 60.2500 381.2000 60.5500 ;
      RECT 0.0000 57.5500 381.2000 60.2500 ;
      RECT 0.6200 57.2500 381.2000 57.5500 ;
      RECT 0.0000 54.5500 381.2000 57.2500 ;
      RECT 0.6200 54.2500 381.2000 54.5500 ;
      RECT 0.0000 51.5500 381.2000 54.2500 ;
      RECT 0.6200 51.2500 381.2000 51.5500 ;
      RECT 0.0000 48.5500 381.2000 51.2500 ;
      RECT 0.6200 48.2500 381.2000 48.5500 ;
      RECT 0.0000 45.5500 381.2000 48.2500 ;
      RECT 0.6200 45.2500 381.2000 45.5500 ;
      RECT 0.0000 42.5500 381.2000 45.2500 ;
      RECT 0.6200 42.2500 381.2000 42.5500 ;
      RECT 0.0000 39.5500 381.2000 42.2500 ;
      RECT 0.6200 39.2500 381.2000 39.5500 ;
      RECT 0.0000 36.5500 381.2000 39.2500 ;
      RECT 0.6200 36.2500 381.2000 36.5500 ;
      RECT 0.0000 33.5500 381.2000 36.2500 ;
      RECT 0.6200 33.2500 381.2000 33.5500 ;
      RECT 0.0000 30.5500 381.2000 33.2500 ;
      RECT 0.6200 30.2500 381.2000 30.5500 ;
      RECT 0.0000 27.5500 381.2000 30.2500 ;
      RECT 0.6200 27.2500 381.2000 27.5500 ;
      RECT 0.0000 24.5500 381.2000 27.2500 ;
      RECT 0.6200 24.2500 381.2000 24.5500 ;
      RECT 0.0000 21.5500 381.2000 24.2500 ;
      RECT 0.6200 21.2500 381.2000 21.5500 ;
      RECT 0.0000 18.5500 381.2000 21.2500 ;
      RECT 0.6200 18.2500 381.2000 18.5500 ;
      RECT 0.0000 15.5500 381.2000 18.2500 ;
      RECT 0.6200 15.2500 381.2000 15.5500 ;
      RECT 0.0000 12.5500 381.2000 15.2500 ;
      RECT 0.6200 12.2500 381.2000 12.5500 ;
      RECT 0.0000 9.5500 381.2000 12.2500 ;
      RECT 0.6200 9.2500 381.2000 9.5500 ;
      RECT 0.0000 6.5500 381.2000 9.2500 ;
      RECT 0.6200 6.2500 381.2000 6.5500 ;
      RECT 0.0000 3.5500 381.2000 6.2500 ;
      RECT 0.6200 3.2500 381.2000 3.5500 ;
      RECT 0.0000 1.3500 381.2000 3.2500 ;
      RECT 0.6200 1.0500 381.2000 1.3500 ;
      RECT 0.0000 0.0000 381.2000 1.0500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 381.2000 380.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 381.2000 380.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 381.2000 380.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 381.2000 380.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 381.2000 380.0000 ;
  END
END core

END LIBRARY
